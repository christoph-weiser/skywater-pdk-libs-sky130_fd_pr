* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param capunits=1.0e-6
.param dkisepp5x=0.745
.param dknfpp=1.0
.param dknfpp5x=1.0009
.param sky130_fd_pr__special_nfet_pass_flash__cdsc_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cdscb_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cdscd_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cit_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__special_nfet_pass_flash__dvt0_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dwg_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_flash__k2_diff_1=0.0
.param sky130_fd_pr__special_nfet_pass_flash__k3_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__kt1_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_flash__kt1l_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__kt2_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__lint_slope=0.0
.param sky130_fd_pr__special_nfet_pass_flash__nfactor_slope=0.0
.param sky130_fd_pr__special_nfet_pass_flash__nlx_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__tox_slope=0.006589
.param sky130_fd_pr__special_nfet_pass_flash__voff_slope=0.0
.param sky130_fd_pr__special_nfet_pass_flash__vth0_slope=0.010889
.param sky130_fd_pr__special_nfet_pass_flash__wint_slope=0.0
.param globalk=1.0
.param hv_dlc_rotweak=0.0
.param localkswitch=1.0
.param lv_dlc_rotweak=0.0
.param lvhvt_dlc_rotweak=0.0
.param lvt_dlc_rotweak=0.0
.param mcl1p1f_cc_w_1_200_s_5_250=0.0
.param mcm1l1d_cc_w_1_360_s_0_360=3.25e-11
.param mcm2d_cc_w_0_140_s_1_540=2.6e-11
.param mcm2m1l1_cc_w_1_120_s_3_500=5.0e-14
.param mcm2p1f_cc_w_1_200_s_0_420=4.11e-11
.param mcm3m2_cc_w_0_300_s_3_300=9.9e-12
.param mcm4m2f_cf_w_1_120_s_0_140=2.69e-12
.param mcm5m1p1_cc_w_0_140_s_0_840=3.22e-11
.param mcm5m2f_cc_w_1_120_s_0_840=4.63e-11
.param mcm5m4_cc_w_1_600_s_10_000=4.0e-12
.param mcm5m4m3_cc_w_2_400_s_9_000=5.0e-14
.param mcrdlm3m2_cc_w_0_300_s_2_100=1.55e-11
.param mcrdlm4l1_cc_w_0_300_s_3_300=1.91e-11
.param mcrdlm4p1_cc_w_0_300_s_3_300=2.02e-11
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ku0_diff=-4.5e-8
.param sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff=0.3
.param sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff=1.1e-8
.param sky130_fd_pr__nfet_g5v0d10v5__lint_slope=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__lku0_diff=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope=0.12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_lint_slope=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope=0.12
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope=0.008
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1=0.0205
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope2=0.01
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope3=0.0067
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope=0.13
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_vth0_slope=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_wint_slope=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__lint1_slope=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__lint_slope=3.0e-9
.param sky130_fd_pr__rf_nfet_g5v0d10v5__nfactor_slope=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox2_slope=0.0086
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox3_slope=0.0055
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox4_slope=0.0255
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox_offset=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__tox_slope=0.008
.param sky130_fd_pr__rf_nfet_g5v0d10v5__voff2_slope=0.0085
.param sky130_fd_pr__rf_nfet_g5v0d10v5__voff_slope=0.00375
.param sky130_fd_pr__rf_nfet_g5v0d10v5__wint_slope=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rshn_mult=1.0
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope=0.008
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1=0.0205
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2=0.01
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3=0.0067
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_slope=0.13
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_slope=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__wint_slope=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__wku0_diff=2.0e-7
.param sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff=6.5e-7
.param sky130_fd_pr__nfet_g5v0d10v5__wlod_diff=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult=1.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ku0_diff=-3.0e-8
.param sky130_fd_pr__nfet_05v0_nvt__kvsat_diff=0.4
.param sky130_fd_pr__nfet_05v0_nvt__kvth0_diff=-7.0e-9
.param sky130_fd_pr__nfet_05v0_nvt__lint_slope=0.0
.param sky130_fd_pr__nfet_05v0_nvt__lku0_diff=0.0
.param sky130_fd_pr__nfet_05v0_nvt__lkvth0_diff=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_slope=0.02
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_05v0_nvt__toxe_slope=0.00105
.param sky130_fd_pr__nfet_05v0_nvt__toxe_slope1=0.01205
.param sky130_fd_pr__nfet_05v0_nvt__toxe_slope2=0.02525
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_slope=0.0035
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_slope=0.0012
.param sky130_fd_pr__nfet_05v0_nvt__wint_slope=0.0
.param sky130_fd_pr__nfet_05v0_nvt__wku0_diff=2.0e-7
.param sky130_fd_pr__nfet_05v0_nvt__wkvth0_diff=8.0e-7
.param sky130_fd_pr__nfet_05v0_nvt__wlod_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak=lvt_dlc_rotweak
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ku0_diff=-2.7e-8
.param sky130_fd_pr__nfet_01v8_lvt__kvsat_diff=0.2
.param sky130_fd_pr__nfet_01v8_lvt__kvth0_diff=7.9e-9
.param sky130_fd_pr__nfet_01v8_lvt__lint_slope=0.0
.param sky130_fd_pr__nfet_01v8_lvt__lku0_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_slope=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__b_toxe_slope=0.003443
.param sky130_fd_pr__rf_nfet_01v8_lvt__b_vth0_slope=0.006056
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__base__dlc_rotweak=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__toxe1_slope=0.008089
.param sky130_fd_pr__rf_nfet_01v8_lvt__toxe_slope=0.006789
.param sky130_fd_pr__nfet_01v8_lvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope=0.003443
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope1=0.002443
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_slope=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope=0.005456
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope1=0.005456
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope2=0.007456
.param sky130_fd_pr__nfet_01v8_lvt__wint_slope=0.0
.param sky130_fd_pr__nfet_01v8_lvt__wku0_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff=3.0e-7
.param sky130_fd_pr__nfet_01v8_lvt__wlod_diff=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__ua_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__ub_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__cdsc_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cdscb_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cdscd_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cit_diff=0.0
.param sky130_fd_pr__special_nfet_pass__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__special_nfet_pass__dvt0_diff=0.0
.param sky130_fd_pr__special_nfet_pass__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__k3_diff=0.0
.param sky130_fd_pr__special_nfet_pass__kt1_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__kt1l_diff=0.0
.param sky130_fd_pr__special_nfet_pass__kt2_diff=0.0
.param sky130_fd_pr__special_nfet_pass__lint_slope=0.0
.param sky130_fd_pr__special_nfet_pass__nfactor_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__nfactor_slope=0.0
.param sky130_fd_pr__special_nfet_pass__rdsw_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__tox_slope=0.003589
.param sky130_fd_pr__special_nfet_pass__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__voff_slope=0.0
.param sky130_fd_pr__special_nfet_pass__vsat_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__vth0_slope=0.005589
.param sky130_fd_pr__special_nfet_pass__wint_slope=0.0
.param sky130_fd_pr__special_nfet_pass_lowleakage__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__special_nfet_latch__cdsc_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cdscb_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cdscd_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cit_diff=0.0
.param sky130_fd_pr__special_nfet_latch__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__special_nfet_latch__dvt0_diff=0.0
.param sky130_fd_pr__special_nfet_latch__dvt1_diff=0.0
.param sky130_fd_pr__special_nfet_latch__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__k3_diff=0.0
.param sky130_fd_pr__special_nfet_latch__kt1_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__kt2_diff=0.0
.param sky130_fd_pr__special_nfet_latch__lint_slope=0.0
.param sky130_fd_pr__special_nfet_latch__nfactor_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__nfactor_slope=0.0
.param sky130_fd_pr__special_nfet_latch__rdsw_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__tox_slope=0.005989
.param sky130_fd_pr__special_nfet_latch__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__voff_slope=0.0
.param sky130_fd_pr__special_nfet_latch__vsat_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__vth0_slope=0.005289
.param sky130_fd_pr__special_nfet_latch__wint_slope=0.0
.param sky130_fd_pr__special_nfet_latch_lowleakage__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__lint_slope=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_slope=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
.param sky130_fd_pr__rf_nfet_01v8__b_toxe_slope=0.003443
.param sky130_fd_pr__rf_nfet_01v8__b_voff_slope=0.007
.param sky130_fd_pr__rf_nfet_01v8__b_vth0_slope=0.005556
.param sky130_fd_pr__rf_nfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8__lint1_slope=0.0
.param sky130_fd_pr__rf_nfet_01v8__lint_slope=5.767e-9
.param sky130_fd_pr__rf_nfet_01v8__toxe1_slope=0.006989
.param sky130_fd_pr__rf_nfet_01v8__toxe2_slope=0.005989
.param sky130_fd_pr__rf_nfet_01v8__toxe3_slope=0.01089
.param sky130_fd_pr__rf_nfet_01v8__toxe4_slope=0.01289
.param sky130_fd_pr__rf_nfet_01v8__toxe_slope=0.008989
.param sky130_fd_pr__nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8__toxe_slope=0.003443
.param sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__voff_slope=0.007
.param sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope=0.003356
.param sky130_fd_pr__nfet_01v8__vth0_slope1=0.007356
.param sky130_fd_pr__nfet_01v8__wint_slope=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ku0_diff=-3.0e-8
.param sky130_fd_pr__nfet_03v3_nvt__kvsat_diff=0.3
.param sky130_fd_pr__nfet_03v3_nvt__kvth0_diff=-2.0e-9
.param sky130_fd_pr__nfet_03v3_nvt__lint_slope=0.0
.param sky130_fd_pr__nfet_03v3_nvt__lku0_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__lkvth0_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_slope=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__toxe_slope=0.0045
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_slope=0.0065
.param sky130_fd_pr__nfet_03v3_nvt__vth0_slope=0.006
.param sky130_fd_pr__nfet_03v3_nvt__wint_slope=0.0
.param sky130_fd_pr__nfet_03v3_nvt__wku0_diff=5.0e-7
.param sky130_fd_pr__nfet_03v3_nvt__wkvth0_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__wlod_diff=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__a0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__a0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__a0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__a0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__a0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__agidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ags_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ags_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ags_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ags_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ags_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b1_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b1_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b1_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b1_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__b1_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__bgidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__cgidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__dsub_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__k2_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__k2_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__k2_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__k2_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__k2_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__keta_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__keta_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__keta_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__keta_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__keta_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__kt2_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ku0_diff=-9.9e-8
.param sky130_fd_pr__nfet_g5v0d16v0__kvsat_diff=0.3
.param sky130_fd_pr__nfet_g5v0d16v0__kvth0_diff=1.7057e-8
.param sky130_fd_pr__nfet_g5v0d16v0__lku0_diff=9.6975e-7
.param sky130_fd_pr__nfet_g5v0d16v0__lkvth0_diff=2.2691e-7
.param sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__nfactor_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ua_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ua_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ua_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ua_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ua_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ub_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ub_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ub_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ub_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ub_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ute_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ute_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ute_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ute_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__ute_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__voff_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__voff_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__voff_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__voff_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__voff_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d16v0__wku0_diff=2.0e-7
.param sky130_fd_pr__nfet_g5v0d16v0__wkvth0_diff=2.3093e-6
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__dlc_rotweak=lvhvt_dlc_rotweak
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__lint_slope=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope=0.005
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope=0.01
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope=0.0055
.param sky130_fd_pr__pfet_01v8_hvt__wint_slope=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ku0_diff=7.0e-8
.param sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff=0.4
.param sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff=3.5e-8
.param sky130_fd_pr__pfet_g5v0d10v5__lint_slope=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__lku0_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope=0.02
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rshp_mult=1.0
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope=0.012
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1=0.02
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2=0.023
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3=0.014
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_slope=0.009
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_slope=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__wint_slope=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__wku0_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff=6.5e-7
.param sky130_fd_pr__pfet_g5v0d10v5__wlod_diff=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult=1.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__dlc_rotweak=lvt_dlc_rotweak
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ku0_diff=5.9e-8
.param sky130_fd_pr__pfet_01v8_lvt__kvsat_diff=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kvth0_diff=1.76e-8
.param sky130_fd_pr__pfet_01v8_lvt__lint_slope=0.0
.param sky130_fd_pr__pfet_01v8_lvt__lku0_diff=0.0
.param sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rf_base_dlc_rotweak=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope=0.003689
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope1=0.01489
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope2=0.01689
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope3=0.02389
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope=0.01389
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope1=0.009789
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope2=0.01089
.param sky130_fd_pr__pfet_01v8_lvt__wint_slope=0.0
.param sky130_fd_pr__pfet_01v8_lvt__wku0_diff=0.0
.param sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff=7.3e-7
.param sky130_fd_pr__pfet_01v8_lvt__wlod_diff=0.0
.param sky130_fd_pr__pfet_01v8_mvt__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__nfactor_slope=0.1
.param sky130_fd_pr__pfet_01v8_mvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_mvt__aw_rd_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_mvt__aw_rs_mult=1.0
.param sky130_fd_pr__pfet_01v8_mvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_mvt__toxe_slope=0.025
.param sky130_fd_pr__pfet_01v8_mvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__ua_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__ua_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__ub_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__ub_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__voff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_mvt__voff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_mvt__voff_slope=0.0
.param sky130_fd_pr__pfet_01v8_mvt__vth0_slope=0.05
.param sky130_fd_pr__special_pfet_pass__cdsc_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cdscb_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cdscd_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cit_diff=0.0
.param sky130_fd_pr__special_pfet_pass__dlc_diff=0.0
.param sky130_fd_pr__special_pfet_pass__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__special_pfet_pass__dvt0_diff=0.0
.param sky130_fd_pr__special_pfet_pass__dwc_diff=0.0
.param sky130_fd_pr__special_pfet_pass__k2_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__k3_diff=0.0
.param sky130_fd_pr__special_pfet_pass__kt1_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__kt1l_diff=0.0
.param sky130_fd_pr__special_pfet_pass__kt2_diff=0.0
.param sky130_fd_pr__special_pfet_pass__lint_diff=0.0
.param sky130_fd_pr__special_pfet_pass__lint_slope=0.0
.param sky130_fd_pr__special_pfet_pass__nfactor_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__nfactor_slope=0.0
.param sky130_fd_pr__special_pfet_pass__rdsw_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__tox_mult=1.0
.param sky130_fd_pr__special_pfet_pass__tox_slope=0.005567
.param sky130_fd_pr__special_pfet_pass__voff_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__voff_slope=0.0
.param sky130_fd_pr__special_pfet_pass__vsat_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__vth0_slope=0.005567
.param sky130_fd_pr__special_pfet_pass__wint_diff=0.0
.param sky130_fd_pr__special_pfet_pass__wint_slope=0.0
.param sky130_fd_pr__special_pfet_pass_lowleakage__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__pfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__dlc_rotweak=lv_dlc_rotweak
.param sky130_fd_pr__pfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ku0_diff=4.5e-8
.param sky130_fd_pr__pfet_01v8__kvsat_diff=0.5
.param sky130_fd_pr__pfet_01v8__kvth0_diff=3.29e-8
.param sky130_fd_pr__pfet_01v8__lint_slope=0.0
.param sky130_fd_pr__pfet_01v8__lku0_diff=0.0
.param sky130_fd_pr__pfet_01v8__lkvth0_diff=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope=0.1
.param sky130_fd_pr__pfet_01v8__nfactor_slope1=0.1
.param sky130_fd_pr__pfet_01v8__nfactor_slope2=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_9=0.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rd_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rs_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1=0.1
.param sky130_fd_pr__rf_pfet_01v8__b_toxe_slope=0.006443
.param sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1=0.004443
.param sky130_fd_pr__rf_pfet_01v8__b_voff_slope=0.014
.param sky130_fd_pr__rf_pfet_01v8__b_voff_slope1=0.009
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1=0.007356
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2=0.009356
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3=0.008356
.param sky130_fd_pr__rf_pfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8__base__dlc_rotweak=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8__nfactor1_slope=0.0
.param sky130_fd_pr__rf_pfet_01v8__nfactor_slope=0.429
.param sky130_fd_pr__rf_pfet_01v8__toxe1_slope=0.01067
.param sky130_fd_pr__rf_pfet_01v8__toxe2_slope=0.01167
.param sky130_fd_pr__rf_pfet_01v8__toxe3_slope=0.01367
.param sky130_fd_pr__rf_pfet_01v8__toxe4_slope=0.01467
.param sky130_fd_pr__rf_pfet_01v8__toxe5_slope=0.01567
.param sky130_fd_pr__rf_pfet_01v8__toxe_slope=0.01267
.param sky130_fd_pr__pfet_01v8__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8__toxe_slope=0.004443
.param sky130_fd_pr__pfet_01v8__toxe_slope1=0.006443
.param sky130_fd_pr__pfet_01v8__toxe_slope2=0.003443
.param sky130_fd_pr__pfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__voff_slope=0.0
.param sky130_fd_pr__pfet_01v8__voff_slope1=0.0
.param sky130_fd_pr__pfet_01v8__voff_slope2=0.007
.param sky130_fd_pr__pfet_01v8__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__vth0_slope=0.005856
.param sky130_fd_pr__pfet_01v8__vth0_slope1=0.007356
.param sky130_fd_pr__pfet_01v8__vth0_slope2=0.004356
.param sky130_fd_pr__pfet_01v8__wint_slope=0.0
.param sky130_fd_pr__pfet_01v8__wku0_diff=2.5e-7
.param sky130_fd_pr__pfet_01v8__wkvth0_diff=2.0e-7
.param sky130_fd_pr__pfet_01v8__wlod_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__a0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__a0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ags_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ags_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbacc_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbacc_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbinv_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbinv_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigc_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigc_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bigsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bigsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cf_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cjswgs_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__pfet_g5v0d16v0__dsub_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__dsub_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__jtssws_diff_0=-4.02e-12
.param sky130_fd_pr__pfet_g5v0d16v0__jtssws_diff_1=-4.02e-12
.param sky130_fd_pr__pfet_g5v0d16v0__k2_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__k2_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__keta_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__keta_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ku0_diff=2.218e-7
.param sky130_fd_pr__pfet_g5v0d16v0__kvsat_diff=0.4
.param sky130_fd_pr__pfet_g5v0d16v0__kvth0_diff=5.2302e-9
.param sky130_fd_pr__pfet_g5v0d16v0__lku0_diff=8.7129e-7
.param sky130_fd_pr__pfet_g5v0d16v0__lkvth0_diff=-4.8631e-7
.param sky130_fd_pr__pfet_g5v0d16v0__lpe0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__lpe0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nigbacc_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nigbacc_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nigbinv_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nigbinv_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rshp_mult=1.0
.param sky130_fd_pr__pfet_g5v0d16v0__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ua_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ua_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ub_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ub_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__voff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__voff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__wku0_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__wkvth0_diff=5.398e-7
.param sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__dlc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_bs_flash__special_sonosfet_star__dwc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__k2_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__k2_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0=-0.44275
.param sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_1=-0.3267
.param sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_2=-0.67944
.param sky130_fd_bs_flash__special_sonosfet_star__lint_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__overlap_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__tox_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope=0.002
.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope1=0.002
.param sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0=-0.0069221
.param sky130_fd_bs_flash__special_sonosfet_star__u0_diff_1=-0.0041919
.param sky130_fd_bs_flash__special_sonosfet_star__u0_diff_2=-0.0081788
.param sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__voff_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__voff_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0=0.91203
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_1=1.3659
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_2=0.27494
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope=0.0255
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope1=0.028
.param sky130_fd_bs_flash__special_sonosfet_star__wint_diff=0.0
.param sonos_eeol_dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_bs_flash__special_sonosfet_original__ajunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__dlc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_bs_flash__special_sonosfet_original__dwc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__k2_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__k2_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__k2_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_0=-0.36466
.param sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_1=-0.029107
.param sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_2=-0.65907
.param sky130_fd_bs_flash__special_sonosfet_original__lint_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_0=-0.23845
.param sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_1=1.3597
.param sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_2=1.0202
.param sky130_fd_bs_flash__special_sonosfet_original__overlap_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__pjunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__tox_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__tox_slope=0.005
.param sky130_fd_bs_flash__special_sonosfet_original__u0_diff_0=-0.004
.param sky130_fd_bs_flash__special_sonosfet_original__u0_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__u0_diff_2=0.0013468
.param sky130_fd_bs_flash__special_sonosfet_original__voff_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__voff_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__voff_diff_2=-0.20912
.param sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_1=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_2=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_0=-1.0278
.param sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_1=-0.85561
.param sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_2=-0.15565
.param sky130_fd_bs_flash__special_sonosfet_original__vth0_slope=0.026
.param sky130_fd_bs_flash__special_sonosfet_original__wint_diff=0.0
.param sonos_peol_dlc_rotweak=hv_dlc_rotweak
.param sky130_fd_pr__nfet_20v0_nvt__reverse_tmax='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt__reverse_vds='-0.01'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vbd_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vbd_2='25.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vbs_1='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vds_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vds_2='25.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vgb_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vgb_2='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vgd_1='sky130_fd_pr__nfet_20v0_nvt__tmax_vds_1'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vgd_2='sky130_fd_pr__nfet_20v0_nvt__tmax_vds_2'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vgs_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt__tmax_vgs_2='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_max='sky130_fd_pr__nfet_20v0_nvt__vbs_max'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_max_1='sky130_fd_pr__nfet_20v0_nvt__vbs_max'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_max_2='sky130_fd_pr__nfet_20v0_nvt__vbs_max'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_min='sky130_fd_pr__nfet_20v0_nvt__vbs_min-sky130_fd_pr__nfet_20v0_nvt__vds_max'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_min_1='sky130_fd_pr__nfet_20v0_nvt__vbs_min-sky130_fd_pr__nfet_20v0_nvt__vds_max_1'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_min_2='sky130_fd_pr__nfet_20v0_nvt__vbs_min-sky130_fd_pr__nfet_20v0_nvt__vds_max_2'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_reversemax='0.501'
.param sky130_fd_pr__nfet_20v0_nvt__vbd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_nvt__vbs_max='0.001'
.param sky130_fd_pr__nfet_20v0_nvt__vbs_max_1='0.001'
.param sky130_fd_pr__nfet_20v0_nvt__vbs_min='-2.501'
.param sky130_fd_pr__nfet_20v0_nvt__vbs_min_1='-2.501'
.param sky130_fd_pr__nfet_20v0_nvt__vds_max='36'
.param sky130_fd_pr__nfet_20v0_nvt__vds_max_1='24.501'
.param sky130_fd_pr__nfet_20v0_nvt__vds_max_2='30.001'
.param sky130_fd_pr__nfet_20v0_nvt__vds_min='-0.001'
.param sky130_fd_pr__nfet_20v0_nvt__vds_min_1='-0.001'
.param sky130_fd_pr__nfet_20v0_nvt__vds_min_2='-0.001'
.param sky130_fd_pr__nfet_20v0_nvt__vgb_max='sky130_fd_pr__nfet_20v0_nvt__vgs_max-sky130_fd_pr__nfet_20v0_nvt__vbs_min'
.param sky130_fd_pr__nfet_20v0_nvt__vgb_max_1='sky130_fd_pr__nfet_20v0_nvt__vgs_max_1-sky130_fd_pr__nfet_20v0_nvt__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_nvt__vgb_max_2='sky130_fd_pr__nfet_20v0_nvt__vgs_max_2-sky130_fd_pr__nfet_20v0_nvt__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_nvt__vgb_min='-1*sky130_fd_pr__nfet_20v0_nvt__vgs_max'
.param sky130_fd_pr__nfet_20v0_nvt__vgb_min_1='0-2.5'
.param sky130_fd_pr__nfet_20v0_nvt__vgb_min_2='0-2.5'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_max='sky130_fd_pr__nfet_20v0_nvt__vgs_max'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_max_1='sky130_fd_pr__nfet_20v0_nvt__vgs_max_1'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_max_2='sky130_fd_pr__nfet_20v0_nvt__vgs_max_2'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_min='-1*sky130_fd_pr__nfet_20v0_nvt__vds_max'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_min_1='-1*sky130_fd_pr__nfet_20v0_nvt__vds_max_1'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_min_2='-1*sky130_fd_pr__nfet_20v0_nvt__vds_max_2'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_reversemax_1='0.101'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_nvt__vgd_reversemin_1='-0.101'
.param sky130_fd_pr__nfet_20v0_nvt__vgs_max='6.501'
.param sky130_fd_pr__nfet_20v0_nvt__vgs_max_1='5.751'
.param sky130_fd_pr__nfet_20v0_nvt__vgs_max_2='6.001'
.param sky130_fd_pr__nfet_20v0_nvt__vgs_min='-1*6.501'
.param sky130_fd_pr__nfet_20v0_nvt__vgs_min_1='-1*5.751'
.param sky130_fd_pr__nfet_20v0_nvt__vgs_min_2='-1*6.001'
.param sky130_fd_pr__nfet_20v0_nvt__vsd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_nvt__vsd_reversemin='-0.501'
.param sky130_fd_pr__nfet_20v0_nvt__vtx='0.020'
.param sky130_fd_pr__nfet_20v0_nvt_iso__k2_diff=-0.11937
.param sky130_fd_pr__nfet_20v0_nvt_iso__reverse_tmax='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__reverse_vds='-0.01'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vbd_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vbd_2='25.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vbs_1='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_2='25.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgb_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgb_2='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgd_1='sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_1'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgd_2='sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vds_2'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgs_1='100.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__tmax_vgs_2='20.001n'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_max='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_max_1='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_max_2='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_min='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min-sky130_fd_pr__nfet_20v0_nvt_iso__vds_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_min_1='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min-sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_min_2='sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min-sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_reversemax='0.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max='0.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbs_max_1='0.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min='-2.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1='-2.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vds_max='22.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1='22.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2='22.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vds_min='-0.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vds_min_1='-0.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vds_min_2='-0.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgb_max='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max-sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgb_max_1='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1-sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgb_max_2='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2-sky130_fd_pr__nfet_20v0_nvt_iso__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgb_min='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgb_min_1='0-2.5'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgb_min_2='0-2.5'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_max='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_max_1='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_max_2='sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_min='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_min_1='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_1'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_min_2='-1*sky130_fd_pr__nfet_20v0_nvt_iso__vds_max_2'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemax_1='0.101'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgd_reversemin_1='-0.101'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max='6.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_1='5.751'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgs_max_2='6.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgs_min='-1*6.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgs_min_1='-1*5.751'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vgs_min_2='-1*6.001'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vsd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vsd_reversemin='-0.501'
.param sky130_fd_pr__nfet_20v0_nvt_iso__vtx='0.02'
.param sky130_fd_pr__nfet_20v0__reverse_tmax='20.001n'
.param sky130_fd_pr__nfet_20v0__reverse_vds='-0.01'
.param sky130_fd_pr__nfet_20v0__rshn_mult=1.0
.param sky130_fd_pr__nfet_20v0__tmax_vbd_1='100.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vbd_2='25.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vbs_1='20.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vds_1='100.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vds_2='25.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vgb_1='100.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vgb_2='20.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vgd_1='sky130_fd_pr__nfet_20v0__tmax_vds_1'
.param sky130_fd_pr__nfet_20v0__tmax_vgd_2='sky130_fd_pr__nfet_20v0__tmax_vds_2'
.param sky130_fd_pr__nfet_20v0__tmax_vgs_1='100.001n'
.param sky130_fd_pr__nfet_20v0__tmax_vgs_2='20.001n'
.param sky130_fd_pr__nfet_20v0__vbd_max='sky130_fd_pr__nfet_20v0__vbs_max'
.param sky130_fd_pr__nfet_20v0__vbd_max_1='sky130_fd_pr__nfet_20v0__vbs_max'
.param sky130_fd_pr__nfet_20v0__vbd_max_2='sky130_fd_pr__nfet_20v0__vbs_max'
.param sky130_fd_pr__nfet_20v0__vbd_min='sky130_fd_pr__nfet_20v0__vbs_min-sky130_fd_pr__nfet_20v0__vds_max'
.param sky130_fd_pr__nfet_20v0__vbd_min_1='sky130_fd_pr__nfet_20v0__vbs_min-sky130_fd_pr__nfet_20v0__vds_max_1'
.param sky130_fd_pr__nfet_20v0__vbd_min_2='sky130_fd_pr__nfet_20v0__vbs_min-sky130_fd_pr__nfet_20v0__vds_max_2'
.param sky130_fd_pr__nfet_20v0__vbd_reversemax='0.501'
.param sky130_fd_pr__nfet_20v0__vbd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0__vbs_max='0.001'
.param sky130_fd_pr__nfet_20v0__vbs_max_1='0.001'
.param sky130_fd_pr__nfet_20v0__vbs_min='-2.501'
.param sky130_fd_pr__nfet_20v0__vbs_min_1='-2.501'
.param sky130_fd_pr__nfet_20v0__vds_max='36'
.param sky130_fd_pr__nfet_20v0__vds_max_1='24.501'
.param sky130_fd_pr__nfet_20v0__vds_max_2='30.001'
.param sky130_fd_pr__nfet_20v0__vds_min='-0.001'
.param sky130_fd_pr__nfet_20v0__vds_min_1='-0.001'
.param sky130_fd_pr__nfet_20v0__vds_min_2='-0.001'
.param sky130_fd_pr__nfet_20v0__vgb_max='sky130_fd_pr__nfet_20v0__vgs_max-sky130_fd_pr__nfet_20v0__vbs_min'
.param sky130_fd_pr__nfet_20v0__vgb_max_1='sky130_fd_pr__nfet_20v0__vgs_max_1-sky130_fd_pr__nfet_20v0__vbs_min_1'
.param sky130_fd_pr__nfet_20v0__vgb_max_2='sky130_fd_pr__nfet_20v0__vgs_max_2-sky130_fd_pr__nfet_20v0__vbs_min_1'
.param sky130_fd_pr__nfet_20v0__vgb_min='-1*sky130_fd_pr__nfet_20v0__vgs_max'
.param sky130_fd_pr__nfet_20v0__vgb_min_1='0-2.5'
.param sky130_fd_pr__nfet_20v0__vgb_min_2='0-2.5'
.param sky130_fd_pr__nfet_20v0__vgd_max='sky130_fd_pr__nfet_20v0__vgs_max'
.param sky130_fd_pr__nfet_20v0__vgd_max_1='sky130_fd_pr__nfet_20v0__vgs_max_1'
.param sky130_fd_pr__nfet_20v0__vgd_max_2='sky130_fd_pr__nfet_20v0__vgs_max_2'
.param sky130_fd_pr__nfet_20v0__vgd_min='-1*sky130_fd_pr__nfet_20v0__vds_max'
.param sky130_fd_pr__nfet_20v0__vgd_min_1='-1*sky130_fd_pr__nfet_20v0__vds_max_1'
.param sky130_fd_pr__nfet_20v0__vgd_min_2='-1*sky130_fd_pr__nfet_20v0__vds_max_2'
.param sky130_fd_pr__nfet_20v0__vgd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0__vgd_reversemax_1='0.101'
.param sky130_fd_pr__nfet_20v0__vgd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0__vgd_reversemin_1='-0.101'
.param sky130_fd_pr__nfet_20v0__vgs_max='6.501'
.param sky130_fd_pr__nfet_20v0__vgs_max_1='5.751'
.param sky130_fd_pr__nfet_20v0__vgs_max_2='6.001'
.param sky130_fd_pr__nfet_20v0__vgs_min='-1*6.501'
.param sky130_fd_pr__nfet_20v0__vgs_min_1='-1*5.751'
.param sky130_fd_pr__nfet_20v0__vgs_min_2='-1*6.001'
.param sky130_fd_pr__nfet_20v0__vsd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0__vsd_reversemin='-0.501'
.param sky130_fd_pr__nfet_20v0__vtx='0.623'
.param sky130_fd_pr__nfet_20v0_iso__reverse_tmax='20.001n'
.param sky130_fd_pr__nfet_20v0_iso__reverse_vds='-0.01'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vbd_1='100.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vbd_2='25.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vbs_1='20.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vds_1='100.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vds_2='25.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vgb_1='100.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vgb_2='20.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vgd_1='sky130_fd_pr__nfet_20v0_iso__tmax_vds_1'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vgd_2='sky130_fd_pr__nfet_20v0_iso__tmax_vds_2'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vgs_1='100.001n'
.param sky130_fd_pr__nfet_20v0_iso__tmax_vgs_2='20.001n'
.param sky130_fd_pr__nfet_20v0_iso__vbd_max='sky130_fd_pr__nfet_20v0_iso__vbs_max'
.param sky130_fd_pr__nfet_20v0_iso__vbd_max_1='sky130_fd_pr__nfet_20v0_iso__vbs_max'
.param sky130_fd_pr__nfet_20v0_iso__vbd_max_2='sky130_fd_pr__nfet_20v0_iso__vbs_max'
.param sky130_fd_pr__nfet_20v0_iso__vbd_min='sky130_fd_pr__nfet_20v0_iso__vbs_min-sky130_fd_pr__nfet_20v0_iso__vds_max'
.param sky130_fd_pr__nfet_20v0_iso__vbd_min_1='sky130_fd_pr__nfet_20v0_iso__vbs_min-sky130_fd_pr__nfet_20v0_iso__vds_max_1'
.param sky130_fd_pr__nfet_20v0_iso__vbd_min_2='sky130_fd_pr__nfet_20v0_iso__vbs_min-sky130_fd_pr__nfet_20v0_iso__vds_max_2'
.param sky130_fd_pr__nfet_20v0_iso__vbd_reversemax='0.501'
.param sky130_fd_pr__nfet_20v0_iso__vbd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_iso__vbs_max='0.001'
.param sky130_fd_pr__nfet_20v0_iso__vbs_max_1='0.001'
.param sky130_fd_pr__nfet_20v0_iso__vbs_min='-2.501'
.param sky130_fd_pr__nfet_20v0_iso__vbs_min_1='-2.501'
.param sky130_fd_pr__nfet_20v0_iso__vds_max='22.501'
.param sky130_fd_pr__nfet_20v0_iso__vds_max_1='22.001'
.param sky130_fd_pr__nfet_20v0_iso__vds_max_2='22.001'
.param sky130_fd_pr__nfet_20v0_iso__vds_min='-0.001'
.param sky130_fd_pr__nfet_20v0_iso__vds_min_1='-0.001'
.param sky130_fd_pr__nfet_20v0_iso__vds_min_2='-0.001'
.param sky130_fd_pr__nfet_20v0_iso__vgb_max='sky130_fd_pr__nfet_20v0_iso__vgs_max-sky130_fd_pr__nfet_20v0_iso__vbs_min'
.param sky130_fd_pr__nfet_20v0_iso__vgb_max_1='sky130_fd_pr__nfet_20v0_iso__vgs_max_1-sky130_fd_pr__nfet_20v0_iso__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_iso__vgb_max_2='sky130_fd_pr__nfet_20v0_iso__vgs_max_2-sky130_fd_pr__nfet_20v0_iso__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_iso__vgb_min='-1*sky130_fd_pr__nfet_20v0_iso__vgs_max'
.param sky130_fd_pr__nfet_20v0_iso__vgb_min_1='0-2.5'
.param sky130_fd_pr__nfet_20v0_iso__vgb_min_2='0-2.5'
.param sky130_fd_pr__nfet_20v0_iso__vgd_max='sky130_fd_pr__nfet_20v0_iso__vgs_max'
.param sky130_fd_pr__nfet_20v0_iso__vgd_max_1='sky130_fd_pr__nfet_20v0_iso__vgs_max_1'
.param sky130_fd_pr__nfet_20v0_iso__vgd_max_2='sky130_fd_pr__nfet_20v0_iso__vgs_max_2'
.param sky130_fd_pr__nfet_20v0_iso__vgd_min='-1*sky130_fd_pr__nfet_20v0_iso__vds_max'
.param sky130_fd_pr__nfet_20v0_iso__vgd_min_1='-1*sky130_fd_pr__nfet_20v0_iso__vds_max_1'
.param sky130_fd_pr__nfet_20v0_iso__vgd_min_2='-1*sky130_fd_pr__nfet_20v0_iso__vds_max_2'
.param sky130_fd_pr__nfet_20v0_iso__vgd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_iso__vgd_reversemax_1='0.101'
.param sky130_fd_pr__nfet_20v0_iso__vgd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_iso__vgd_reversemin_1='-0.101'
.param sky130_fd_pr__nfet_20v0_iso__vgs_max='6.501'
.param sky130_fd_pr__nfet_20v0_iso__vgs_max_1='5.751'
.param sky130_fd_pr__nfet_20v0_iso__vgs_max_2='6.001'
.param sky130_fd_pr__nfet_20v0_iso__vgs_min='-1*6.501'
.param sky130_fd_pr__nfet_20v0_iso__vgs_min_1='-1*5.751'
.param sky130_fd_pr__nfet_20v0_iso__vgs_min_2='-1*6.001'
.param sky130_fd_pr__nfet_20v0_iso__vsd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_iso__vsd_reversemin='-0.501'
.param sky130_fd_pr__nfet_20v0_iso__vtx='0.617'
.param sky130_fd_pr__nfet_20v0_zvt__hvvsat_mult=1.0
.param sky130_fd_pr__nfet_20v0_zvt__k2_diff=0.0
.param sky130_fd_pr__nfet_20v0_zvt__lint_diff=0.0
.param sky130_fd_pr__nfet_20v0_zvt__reverse_tmax='20.001n'
.param sky130_fd_pr__nfet_20v0_zvt__reverse_vds='-0.01'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vbd_1='100.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vbd_2='25.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vbs_1='20.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vds_1='100.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vds_2='25.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgb_1='100.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgb_2='20.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgd_1='sky130_fd_pr__nfet_20v0_zvt__tmax_vds_1'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgd_2='sky130_fd_pr__nfet_20v0_zvt__tmax_vds_2'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgs_1='100.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgs_2='20.001n'
.param sky130_fd_pr__nfet_20v0_zvt__tmax_vgs_model01='0.001n'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_max='sky130_fd_pr__nfet_20v0_zvt__vbs_max'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_max_1='sky130_fd_pr__nfet_20v0_zvt__vbs_max'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_max_2='sky130_fd_pr__nfet_20v0_zvt__vbs_max'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_min='sky130_fd_pr__nfet_20v0_zvt__vbs_min-sky130_fd_pr__nfet_20v0_zvt__vds_max'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_min_1='sky130_fd_pr__nfet_20v0_zvt__vbs_min-sky130_fd_pr__nfet_20v0_zvt__vds_max_1'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_min_2='sky130_fd_pr__nfet_20v0_zvt__vbs_min-sky130_fd_pr__nfet_20v0_zvt__vds_max_2'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_reversemax='0.501'
.param sky130_fd_pr__nfet_20v0_zvt__vbd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_zvt__vbs_max='0.001'
.param sky130_fd_pr__nfet_20v0_zvt__vbs_max_1='0.001'
.param sky130_fd_pr__nfet_20v0_zvt__vbs_min='-2.501'
.param sky130_fd_pr__nfet_20v0_zvt__vbs_min_1='-2.501'
.param sky130_fd_pr__nfet_20v0_zvt__vds_max='30.001'
.param sky130_fd_pr__nfet_20v0_zvt__vds_max_1='24.501'
.param sky130_fd_pr__nfet_20v0_zvt__vds_max_2='28.001'
.param sky130_fd_pr__nfet_20v0_zvt__vds_max_model01='1*3.0'
.param sky130_fd_pr__nfet_20v0_zvt__vds_min='-0.001'
.param sky130_fd_pr__nfet_20v0_zvt__vds_min_1='-0.001'
.param sky130_fd_pr__nfet_20v0_zvt__vds_min_2='-0.001'
.param sky130_fd_pr__nfet_20v0_zvt__vds_min_model01='-1*3.0'
.param sky130_fd_pr__nfet_20v0_zvt__vgb_max='sky130_fd_pr__nfet_20v0_zvt__vgs_max-sky130_fd_pr__nfet_20v0_zvt__vbs_min'
.param sky130_fd_pr__nfet_20v0_zvt__vgb_max_1='sky130_fd_pr__nfet_20v0_zvt__vgs_max_1-sky130_fd_pr__nfet_20v0_zvt__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_zvt__vgb_max_2='sky130_fd_pr__nfet_20v0_zvt__vgs_max_2-sky130_fd_pr__nfet_20v0_zvt__vbs_min_1'
.param sky130_fd_pr__nfet_20v0_zvt__vgb_min='-1*sky130_fd_pr__nfet_20v0_zvt__vgs_max'
.param sky130_fd_pr__nfet_20v0_zvt__vgb_min_1='0-2.5'
.param sky130_fd_pr__nfet_20v0_zvt__vgb_min_2='0-2.5'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_max='sky130_fd_pr__nfet_20v0_zvt__vgs_max'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_max_1='sky130_fd_pr__nfet_20v0_zvt__vgs_max_1'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_max_2='sky130_fd_pr__nfet_20v0_zvt__vgs_max_2'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_min='-1*sky130_fd_pr__nfet_20v0_zvt__vds_max'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_min_1='-1*sky130_fd_pr__nfet_20v0_zvt__vds_max_1'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_min_2='-1*sky130_fd_pr__nfet_20v0_zvt__vds_max_2'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_reversemax_1='0.101'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_reversemin='-5.501'
.param sky130_fd_pr__nfet_20v0_zvt__vgd_reversemin_1='-0.101'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_max='6.501'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_max_1='5.751'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_max_2='6.001'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_max_model01='1*3.0'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_min='-1*6.501'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_min_1='-1*5.751'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_min_2='-1*6.001'
.param sky130_fd_pr__nfet_20v0_zvt__vgs_min_model01='-1*3.0'
.param sky130_fd_pr__nfet_20v0_zvt__vsat_diff=0.0
.param sky130_fd_pr__nfet_20v0_zvt__vsd_reversemax='5.501'
.param sky130_fd_pr__nfet_20v0_zvt__vsd_reversemin='-0.501'
.param sky130_fd_pr__nfet_20v0_zvt__vtx='-0.223'
.param sky130_fd_pr__pfet_20v0__agidl_diff=0.0
.param sky130_fd_pr__pfet_20v0__k2_diff=0.0
.param sky130_fd_pr__pfet_20v0__reverse_tmax='20.001n'
.param sky130_fd_pr__pfet_20v0__reverse_vds='0.01'
.param sky130_fd_pr__pfet_20v0__rshn_mult=1.0
.param sky130_fd_pr__pfet_20v0__tmax_vbd_1='100.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vbd_2='25.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vbs_1='20.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vds_1='100.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vds_2='25.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vgb_1='100.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vgb_2='20.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vgd_1='sky130_fd_pr__pfet_20v0__tmax_vds_1'
.param sky130_fd_pr__pfet_20v0__tmax_vgd_2='sky130_fd_pr__pfet_20v0__tmax_vds_2'
.param sky130_fd_pr__pfet_20v0__tmax_vgs_1='100.001n'
.param sky130_fd_pr__pfet_20v0__tmax_vgs_2='20.001n'
.param sky130_fd_pr__pfet_20v0__vbd_max='sky130_fd_pr__pfet_20v0__vbs_max-sky130_fd_pr__pfet_20v0__vds_min'
.param sky130_fd_pr__pfet_20v0__vbd_max_1='sky130_fd_pr__pfet_20v0__vbs_max-sky130_fd_pr__pfet_20v0__vds_min_1'
.param sky130_fd_pr__pfet_20v0__vbd_max_2='sky130_fd_pr__pfet_20v0__vbs_max-sky130_fd_pr__pfet_20v0__vds_min_2'
.param sky130_fd_pr__pfet_20v0__vbd_min='sky130_fd_pr__pfet_20v0__vbs_min'
.param sky130_fd_pr__pfet_20v0__vbd_min_1='sky130_fd_pr__pfet_20v0__vbs_min'
.param sky130_fd_pr__pfet_20v0__vbd_min_2='sky130_fd_pr__pfet_20v0__vbs_min'
.param sky130_fd_pr__pfet_20v0__vbd_reversemax='5.501'
.param sky130_fd_pr__pfet_20v0__vbd_reversemin='-0.501'
.param sky130_fd_pr__pfet_20v0__vbs_max='2.501'
.param sky130_fd_pr__pfet_20v0__vbs_max_1='2.501'
.param sky130_fd_pr__pfet_20v0__vbs_min='-0.001'
.param sky130_fd_pr__pfet_20v0__vbs_min_1='-0.001'
.param sky130_fd_pr__pfet_20v0__vds_max='0.01'
.param sky130_fd_pr__pfet_20v0__vds_max_1='0.01'
.param sky130_fd_pr__pfet_20v0__vds_max_2='0.01'
.param sky130_fd_pr__pfet_20v0__vds_min='-28.001'
.param sky130_fd_pr__pfet_20v0__vds_min_1='-24.501'
.param sky130_fd_pr__pfet_20v0__vds_min_2='-24.501'
.param sky130_fd_pr__pfet_20v0__vgb_max='-1*sky130_fd_pr__pfet_20v0__vgs_min'
.param sky130_fd_pr__pfet_20v0__vgb_max_1='0+1.0'
.param sky130_fd_pr__pfet_20v0__vgb_max_2='0+1.0'
.param sky130_fd_pr__pfet_20v0__vgb_min='sky130_fd_pr__pfet_20v0__vgs_min-sky130_fd_pr__pfet_20v0__vbs_max'
.param sky130_fd_pr__pfet_20v0__vgb_min_1='sky130_fd_pr__pfet_20v0__vgs_min_1-sky130_fd_pr__pfet_20v0__vbs_max_1'
.param sky130_fd_pr__pfet_20v0__vgb_min_2='sky130_fd_pr__pfet_20v0__vgs_min_2-sky130_fd_pr__pfet_20v0__vbs_max_1'
.param sky130_fd_pr__pfet_20v0__vgd_max='-1*sky130_fd_pr__pfet_20v0__vds_min'
.param sky130_fd_pr__pfet_20v0__vgd_max_1='-1*sky130_fd_pr__pfet_20v0__vds_min_1'
.param sky130_fd_pr__pfet_20v0__vgd_max_2='-1*sky130_fd_pr__pfet_20v0__vds_min_2'
.param sky130_fd_pr__pfet_20v0__vgd_min='sky130_fd_pr__pfet_20v0__vgs_min'
.param sky130_fd_pr__pfet_20v0__vgd_min_1='sky130_fd_pr__pfet_20v0__vgs_min_1'
.param sky130_fd_pr__pfet_20v0__vgd_min_2='sky130_fd_pr__pfet_20v0__vgs_min_2'
.param sky130_fd_pr__pfet_20v0__vgd_reversemax='5.501'
.param sky130_fd_pr__pfet_20v0__vgd_reversemax_1='0.101'
.param sky130_fd_pr__pfet_20v0__vgd_reversemin='-5.501'
.param sky130_fd_pr__pfet_20v0__vgd_reversemin_1='-0.101'
.param sky130_fd_pr__pfet_20v0__vgs_max='-1*-6.501'
.param sky130_fd_pr__pfet_20v0__vgs_max_1='-1*-5.751'
.param sky130_fd_pr__pfet_20v0__vgs_max_2='-1*-6.001'
.param sky130_fd_pr__pfet_20v0__vgs_min='-6.501'
.param sky130_fd_pr__pfet_20v0__vgs_min_1='-5.751'
.param sky130_fd_pr__pfet_20v0__vgs_min_2='-6.001'
.param sky130_fd_pr__pfet_20v0__vsd_reversemax='0.501'
.param sky130_fd_pr__pfet_20v0__vsd_reversemin='-5.501'
.param sky130_fd_pr__pfet_20v0__vtx='-0.873'