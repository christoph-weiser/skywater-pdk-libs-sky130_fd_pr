* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

x0 dw_n700_n714# a_n900_n1000# a_1050_0# subs sky130_fd_pr__nfet_20v0 w=3e+07u l=1.5e+06u
x1 dw_n700_n714# a_n900_n1000# a_n958_0# subs sky130_fd_pr__nfet_20v0 w=3e+07u l=1.5e+06u