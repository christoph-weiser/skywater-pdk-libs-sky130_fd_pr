* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope=3.189e-03
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope1=1.589e-02
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope2=1.789e-02
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope3=2.389e-02
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope=1.2789e-02
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope1=9.2789e-03
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope2=1.0789e-02
.param sky130_fd_pr__pfet_01v8_lvt__lint_slope=0
.param sky130_fd_pr__pfet_01v8_lvt__wint_slope=0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope=0.017