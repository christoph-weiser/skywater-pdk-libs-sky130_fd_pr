* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__esd_nfet_01v8__toxe_mult=1.0
.param sky130_fd_pr__esd_nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__esd_nfet_01v8__overlap_mult=0.9842
.param sky130_fd_pr__esd_nfet_01v8__ajunction_mult=0.99543
.param sky130_fd_pr__esd_nfet_01v8__pjunction_mult=1.0204
.param sky130_fd_pr__esd_nfet_01v8__lint_diff=0.0
.param sky130_fd_pr__esd_nfet_01v8__wint_diff=0.0
.param sky130_fd_pr__esd_nfet_01v8__dlc_diff=-.61491e-9
.param sky130_fd_pr__esd_nfet_01v8__dwc_diff=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_0=3.4854e-11
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_0=-0.00095204
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_0=-0.05413
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_0=0.017628
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_0=-3.6155e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_0=0.0024163
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_0=-0.003544
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_0=-1486.8
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_0=0.33028
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_1=2.339e-11
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_1=-0.00072437
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_1=-0.041786
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_1=-0.0030404
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_1=-1.2496e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_1=-0.0045709
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_1=-0.0029246
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_1=2103.9
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_1=0.2532
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_2=2.8715e-11
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_2=-0.001174
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_2=-0.073442
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_2=0.0032898
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_2=-4.8763e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_2=-0.0047856
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_2=-0.0040656
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_2=3719.6
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_2=0.40322
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_2=0.0
.include "sky130_fd_pr__esd_nfet_01v8.pm3.spice"