* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=1.042
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=1.2
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=0.99758
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=1.1193
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=1.1801
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=-1.21275e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=2.252e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=7.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=-1.21275e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=4.504e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_0=0.037892
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_0=-7490.2
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_0=0.0061192
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_0=-0.0068374
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_1=0.042869
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_1=-5260.5
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_1=0.0082977
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_1=-0.0034898
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_0=-7602.3
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_0=0.028278
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_0=0.0058947
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_0=-0.0070921
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_1=-7404.4
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_1=0.035525
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_1=0.0078725
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_1=-0.0038822
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_2=-8487.7
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_2=0.039934
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_2=0.0052827
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_2=-0.0061567
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_0=0.0053572
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_0=-0.0056999
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_0=0.037862
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_0=86.018
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_1=0.001022
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_1=-0.0060669
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_1=0.032656
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_1=-8977.1
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_2=0.0043107
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_2=-0.011734
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_2=0.025004
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_2=-884.49
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"