* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__esd_nfet_01v8__toxe_mult=1.052
.param sky130_fd_pr__esd_nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__esd_nfet_01v8__overlap_mult=1.0257
.param sky130_fd_pr__esd_nfet_01v8__ajunction_mult=1.2169e+0
.param sky130_fd_pr__esd_nfet_01v8__pjunction_mult=1.2474e+0
.param sky130_fd_pr__esd_nfet_01v8__lint_diff=-1.7325e-8
.param sky130_fd_pr__esd_nfet_01v8__wint_diff=3.2175e-8
.param sky130_fd_pr__esd_nfet_01v8__dlc_diff=-14.422e-9
.param sky130_fd_pr__esd_nfet_01v8__dwc_diff=3.2175e-8
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_0=1.3831e-10
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_0=0.0017582
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_0=-7.8945e-20
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_0=0.062077
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_0=0.0024646
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_0=29832.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_0=0.3284
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_1=1.1282e-10
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_1=-0.017137
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_1=2.3412e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_1=0.055271
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_1=0.0037507
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_1=15696.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_1=-0.27022
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_2=1.2882e-10
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_2=-0.0077745
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_2=-2.6082e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_2=0.056219
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_2=0.0018148
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_2=26605.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_2=-0.44799
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_2=0.0
.include "sky130_fd_pr__esd_nfet_01v8.pm3.spice"