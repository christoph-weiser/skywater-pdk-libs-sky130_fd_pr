* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param cnwvc=0.0
.param diff_cd=0.0
.param hvn_bodyeffect=0.0
.param hvn_diode=0.0
.param hvn_mobility=0.0
.param hvn_saturation=0.0
.param hvn_subvt=0.0
.param hvn_threshold=0.0
.param hvp_bodyeffect=0.0
.param hvp_diode=0.0
.param hvp_mobility=0.0
.param hvp_saturation=0.0
.param hvp_subvt=0.0
.param hvp_threshold=0.0
.param hvtox=0.0
.param ic_cap=0.0
.param ic_res=0.0
.param ic_res_ndiff=0.0
.param ic_res_pdiff=0.0
.param ic_res_poly=0.0
.param ic_res_pwell=0.0
.param lvhp_bodyeffect=0.0
.param lvhp_mobility=0.0
.param lvhp_saturation=0.0
.param lvhp_threshold=0.0
.param lvln_bodyeffect=0.0
.param lvln_mobility=0.0
.param lvln_saturation=0.0
.param lvln_threshold=0.0
.param lvlp_bodyeffect=0.0
.param lvlp_mobility=0.0
.param lvlp_saturation=0.0
.param lvlp_threshold=0.0
.param lvn_bodyeffect=0.0
.param lvn_diode=0.0
.param lvn_mobility=0.0
.param lvn_saturation=0.0
.param lvn_subvt=0.0
.param lvn_threshold=0.0
.param lvp_bodyeffect=0.0
.param lvp_diode=0.0
.param lvp_mobility=0.0
.param lvp_saturation=0.0
.param lvp_subvt=0.0
.param lvp_threshold=0.0
.param lvtox=0.0
.param mim=0.0
.param hvntvn_threshold=0.0
.param sky130_fd_pr__nfet_20v0_nvt=0.0
.param sky130_fd_pr__nfet_20v0_nvt_iso=0.0
.param sky130_fd_pr__nfet_20v0=0.0
.param sky130_fd_pr__nfet_20v0_iso=0.0
.param n20zvtvh1defet=0.0
.param sky130_fd_pr__nfet_20v0_zvt=0.0
.param ndiff_cd=0.0
.param sky130_fd_pr__pfet_20v0=0.0
.param pdiff_cd=0.0
.param sky130_fd_pr__nfet_01v8_lvt=0.0
.param sky130_fd_pr__special_nfet_pass_lvt=0.0
.param sky130_fd_pr__npn_05v5_all=0.0
.param sky130_fd_pr__nfet_g5v0d16v0=0.0
.param sky130_fd_pr__pfet_01v8_mvt=0.0
.param sky130_fd_pr__pnp_05v5_w0p68l0p68=0.0
.param poly_cd=0.0
.param sky130_fd_pr__pfet_01v8=0.0
.param sky130_fd_pr__pfet_g5v0d16v0=0.0
.param well_diode=0.0