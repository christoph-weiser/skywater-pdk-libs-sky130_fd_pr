* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__esd_pfet_g5v0d10v5__toxe_mult=1.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rshp_mult=1.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__overlap_mult=1.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ajunction_mult=1.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pjunction_mult=1.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__lint_diff=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__wint_diff=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__dlc_diff=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__dwc_diff=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_5=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ub_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ags_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__a0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__k2_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__u0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vth0_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__ua_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__nfactor_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__esd_pfet_g5v0d10v5__b1_diff_7=0.0
.include "sky130_fd_pr__esd_pfet_g5v0d10v5.pm3.spice"