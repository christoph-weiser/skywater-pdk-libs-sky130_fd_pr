* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_bs_flash__special_sonosfet_original__tox_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__ajunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__pjunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__overlap_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_original__lint_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__wint_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__dlc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__dwc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__rdsw_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__vth0_diff_0=-1.0887
.param sky130_fd_bs_flash__special_sonosfet_original__u0_diff_0=-4.4130e-3
.param sky130_fd_bs_flash__special_sonosfet_original__vsat_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__voff_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__k2_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_original__nfactor_diff_0=-5.9464e-1
.param sky130_fd_bs_flash__special_sonosfet_original__kt1_diff_0=-3.7039e-1