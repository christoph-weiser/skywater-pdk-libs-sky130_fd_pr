* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult=1.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult=1.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult=0.89805
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult=0.99505
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult=1.0144
.param sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0=0.04749
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0=0.010406
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0=0.001245
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0=0.011822
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0=-3.1273e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0=-1672.2
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0=2.4153e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0=-8.8395e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1=0.044
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1=0.010327
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1=0.0029959
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1=0.013091
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1=-3.0744e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1=-1443.7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1=3.4221e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1=-2.42e-11
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2=0.042379
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2=0.010304
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2=0.0012741
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2=0.012354
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2=-3.1062e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2=-43.451
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2=3.291e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2=-7.333e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3=-1.7201e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3=0.043088
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3=0.010034
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3=0.0010628
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3=0.012223
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3=-3.1021e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3=33.54
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3=3.183e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4=2.7249e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4=-7.6527e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4=0.044539
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4=0.0099796
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4=0.0013927
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4=0.010605
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4=-3.1814e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4=-907.07
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5=-6.1783e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5=8.2128e-11
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5=-0.305
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5=-0.021325
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5=-0.26694
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5=0.047533
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5=-0.0063931
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5=0.009901
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5=-2.089e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6=6.0666e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6=-7.0128e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6=0.045318
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6=0.010019
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6=0.0016874
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6=0.010474
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6=-3.1807e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6=1500.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7=-3.6086e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7=3019.2
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7=9.7977e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7=3.2228e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7=0.06372
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7=0.010207
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7=0.0014468
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7=0.011095
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8=-0.0088519
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8=-0.00064109
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8=-2.2058e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8=-6.7671e-19
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8=5.5348e-11
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8=-0.175
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8=0.0071088
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8=0.0024548
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8=0.010977
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9=0.0014488
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9=0.0037985
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9=0.002075
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9=-3.5584e-7
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9=-191.5
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9=1.3051e-18
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9=-1.3283e-11
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9=0.061417
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10=-0.17848
.param sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10=2.8803e-12
.param sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10=-2502.2
.param sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10=8.2506e-20
.param sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10=0.0031768
.param sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10=0.15934
.param sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10=-0.00045045
.param sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10=0.013013
.param sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10=0.0
.include "sky130_fd_pr__esd_nfet_g5v0d10v5.pm3.spice"