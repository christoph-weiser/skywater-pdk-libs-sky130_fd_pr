* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_lvt__toxe_mult=0.9635
.param sky130_fd_pr__pfet_01v8_lvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_lvt__overlap_mult=0.724
.param sky130_fd_pr__pfet_01v8_lvt__ajunction_mult=9.3001e-1
.param sky130_fd_pr__pfet_01v8_lvt__pjunction_mult=9.3439e-1
.param sky130_fd_pr__pfet_01v8_lvt__lint_diff=1.21275e-8
.param sky130_fd_pr__pfet_01v8_lvt__wint_diff=-2.252e-8
.param sky130_fd_pr__pfet_01v8_lvt__dlc_diff=2.0382e-8
.param sky130_fd_pr__pfet_01v8_lvt__dwc_diff=-2.252e-8
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_0=1.8236e-5
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_0=0.057962
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0=0.04699
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_0=0.1188
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_0=0.051281
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_1=0.030016
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_1=6.3753e-5
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_1=0.053089
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1=0.062335
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_1=0.11351
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_2=0.14251
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_2=0.034025
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_2=-2.9718e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_2=-0.042558
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2=0.068905
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_3=0.12793
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_3=0.033467
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_3=5.3522e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_3=-0.0034386
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3=0.060803
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4=0.035185
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_4=-5.7776e-9
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_4=0.039388
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_4=-0.00015853
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4=2649.7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_4=2.0438e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5=0.1099
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_5=1.6482e-7
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_5=0.036896
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_5=-0.00012951
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5=-24859.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_5=3.3037e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_6=0.19249
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6=0.041047
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_6=0.04499
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_6=0.028443
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_6=-0.00026304
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_7=0.15046
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7=0.033761
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_7=0.085016
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_7=0.04862
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_7=-0.00010679
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_8=0.13976
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8=0.080847
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_8=0.067986
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_8=0.035894
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_8=-0.0003169
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_9=0.13129
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9=0.073616
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_9=0.080573
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_9=0.03877
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_9=-0.00030083
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_10=-0.00028535
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10=0.080406
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_10=0.03088
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_10=0.074414
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_10=0.092733
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_11=-0.00036855
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11=6238.9
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11=0.040634
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_11=0.04248
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_12=0.022657
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_12=0.087754
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_12=-0.00033122
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12=-13671.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12=0.052081
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_12=-5.7847e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_13=0.034147
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_13=-0.0039669
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_13=0.10427
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_13=-0.00021283
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13=0.06929
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_14=0.03164
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_14=-0.012
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_14=0.12605
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_14=-0.00010143
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14=0.044427
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_15=0.040581
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_15=0.0080084
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_15=0.11206
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_15=-0.00027917
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15=0.090708
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_16=0.041067
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_16=0.039408
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_16=0.1007
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_16=-0.00021219
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16=0.078926
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_17=0.034165
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_17=0.055625
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_17=0.097238
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_17=-0.0002235
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17=0.079729
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_18=0.035023
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_18=-0.00012027
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18=-9547.2
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18=0.019246
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_19=-2.3922e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_19=0.02131
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_19=0.091925
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_19=-0.00016727
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19=-18404.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19=0.032189
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_20=0.022835
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_20=0.10505
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_20=0.092125
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_20=-0.00015806
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20=0.042628
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_21=-0.00015959
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21=0.038854
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_21=0.040801
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_21=0.090482
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_21=0.10086
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_22=0.16358
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_22=0.077614
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_22=-0.00011519
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22=0.04077
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_22=1.3e-12
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_22=0.044326
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_23=0.035049
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_23=0.0040365
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_23=0.11133
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_23=-0.00016106
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23=0.072293
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_24=0.032947
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_24=0.022112
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_24=0.11166
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_24=-0.00013292
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24=0.066105
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_25=0.032376
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_25=-0.00010893
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25=2460.8
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25=-0.004201
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_26=0.02304
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_26=0.086586
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_26=-0.00014865
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26=-7093.1
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26=0.030421
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_26=-3.0509e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_27=5.4132e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_27=4.7258e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_27=0.044406
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_27=0.00040064
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27=0.015981
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_28=-6.2589e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_28=2.1373e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_28=0.013052
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_28=-9.9946e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28=0.04864
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_29=1.1353e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_29=2.324e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_29=0.023227
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_29=-3.4446e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29=0.075546
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_30=-2.424e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_30=2.2494e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_30=0.026211
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_30=-4.4666e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30=0.049375
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_31=5.9189e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_31=2.2715e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_31=0.028872
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_31=-0.00012571
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31=0.088628
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_32=6.2247e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32=-5767.1
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32=0.11275
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_32=0.045505
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_33=-6.6705e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33=-19424.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33=0.059647
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_33=1.6932e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_33=2.1062e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_33=0.026212
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_34=0.048415
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_34=-8.0517e-6
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34=0.089735
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_34=1.2734e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_34=3.9757e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_35=0.043931
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_35=-1.3776e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35=0.067319
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_35=5.6032e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_35=1.9598e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_36=0.047583
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_36=-4.5337e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36=0.06697
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_36=9.857e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_36=1.98e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_37=2.1613e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_37=0.034954
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_37=-8.6545e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37=0.057766
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_37=5.8275e-8
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_38=0.032381
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_38=0.00013127
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38=-394.79
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38=-0.014067
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_39=7.5746e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_39=3.4088e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_39=0.021853
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_39=0.00018882
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39=-21675.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39=0.00071188
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_39=0.0
.include "sky130_fd_pr__pfet_01v8_lvt.pm3.spice"