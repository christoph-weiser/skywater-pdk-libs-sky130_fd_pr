* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=0.94
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=0.8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=0.76246
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=0.81753
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=0.77786
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=1.7325e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=-3.2175e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=-7.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=-6.425e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=1.7325e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_0=-0.096862
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_0=-0.33307
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_0=-12674.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_0=-0.0035704
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_0=-0.32676
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_0=-0.0051274
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_1=-0.073057
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_1=-0.50082
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_1=-6173.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_1=-0.011741
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_1=-0.32836
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_1=-0.0039209
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_0=-0.37193
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_0=-12970.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_0=-0.10565
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_0=-0.0039729
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_0=-0.0051626
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_0=-0.28517
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_1=-0.38675
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_1=-8042.9
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_1=-0.080494
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_1=-0.011251
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_1=-0.0041751
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_1=-0.28285
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_2=-0.509
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_2=-9472.9
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_2=-0.082655
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_2=-0.0094809
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_2=-0.0051933
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_2=-0.28355
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_0=-0.0041159
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_0=-0.22789
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_0=-0.0035707
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_0=-0.53245
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_0=-0.096572
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_0=-10255.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_1=-0.016447
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_1=-0.25497
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_1=-0.0053074
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_1=-0.58953
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_1=-0.083034
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_1=-10453.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_2=-0.0084536
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_2=-0.24814
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_2=-0.0025043
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_2=-0.51293
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_2=-0.095613
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_2=-15629.0
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"