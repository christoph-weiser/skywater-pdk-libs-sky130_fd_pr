* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.model sky130_fd_pr__model__parasitic__diode_ps2dn d level=3.0 tlevc=1.0 area=1.0e+12 cj='7.8544e-005*1e-12*sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult' mj=0.49 pb=0.5348 cjsw='8.1664e-010*1e-6*sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult' mjsw=0.20024 php=0.5348 cta=0.0016157 ctp=0.0008 tpb=0.0025003 tphp=0.001675 js=6.1049e-017 jsw=8.1115e-016 n=1.0791 rs=900 ik='2.08e-009/1e-12' ikr='0/1e-12' vb=16.95 ibv=0.00106 trs=0 eg=1.17 xti=1.0 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0