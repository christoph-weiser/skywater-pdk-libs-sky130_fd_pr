* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_g5v0d10v5__toxe_mult=1.0
.param sky130_fd_pr__pfet_g5v0d10v5__rshp_mult=1.0
.param sky130_fd_pr__pfet_g5v0d10v5__overlap_mult=9.8210e-1
.param sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult=1.0050e+0
.param sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult=1.0090e+0
.param sky130_fd_pr__pfet_g5v0d10v5__lint_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__wint_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__dlc_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__dwc_diff=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0=-3.5458e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0=-5.8022e-14
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0=0.014703
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0=0.57788
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0=-0.0014124
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0=-0.028371
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0=-3186.1
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1=-3.0352e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1=6.7649e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1=-0.022679
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1=0.013083
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1=0.283
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1=-0.0014011
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1=-0.021883
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1=-0.042028
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2=-3.6729e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2=3.2719e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2=0.014151
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2=0.50184
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2=-0.0015791
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2=-0.027332
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2=-3569.8
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3=0.001691
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3=-2.6615e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3=-6.9785e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3=0.00019928
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3=0.0057365
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3=0.3885
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3=-0.0007055
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3=-0.0098902
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4=0.46599
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4=-0.00054912
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4=-0.02036
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4=5.3823e-5
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4=-2.8884e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4=-1.2153e-12
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4=0.001753
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4=0.0046061
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5=0.006736
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5=0.54386
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5=-0.0015051
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5=-0.012652
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5=0.013907
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5=-5.0605e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5=-8.9211e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5=-0.0011717
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6=0.011193
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6=0.28744
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6=-0.001941
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6=-0.0018982
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6=-4014.6
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6=-9.2003e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6=-3.2377e-12
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7=0.00058676
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7=0.0089159
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7=-0.011744
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7=0.33401
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7=-0.00081258
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7=-3.1757e-5
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7=-2.5975e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7=-7.3663e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8=-0.022709
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8=0.0071665
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8=-0.0081142
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8=0.39
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8=-0.0010873
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8=-0.039506
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8=-3.9251e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8=-9.5728e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9=0.001555
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9=0.0035952
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9=-0.020147
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9=0.66771
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9=-0.00064541
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9=0.0013478
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9=-1.5597e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9=-4.1075e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10=0.65079
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10=-0.00058739
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10=-0.011509
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10=0.004764
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10=0.0047543
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10=-2.6268e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10=-9.3197e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10=0.00077535
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11=-2669.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11=0.35952
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11=-0.00039781
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11=-0.052985
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11=0.01005
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11=1.6198e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11=-7.89e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12=-2876.4
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12=0.2147
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12=-0.0019672
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12=-0.0056806
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12=0.0064154
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12=-1.3729e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12=-6.0972e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13=-4.7024e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13=-1102.1
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13=0.084251
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13=-0.0010482
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13=-0.036736
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13=0.010768
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13=8.1074e-12
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14=1.4457e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14=-2.7278e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14=-0.022429
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14=0.25329
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14=-0.0012149
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14=-0.025748
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14=-0.043471
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14=0.012945
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15=0.01425
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15=1.0089e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15=-3.7504e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15=-4033.1
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15=0.46809
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15=-0.0015963
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15=-0.030898
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16=-0.01328
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16=-0.019138
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16=0.011784
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16=-7.4832e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16=-6.4597e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16=-0.0087926
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16=0.36309
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16=-0.002041
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17=-0.035514
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17=-0.00037808
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17=-0.02415
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17=0.00030259
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17=0.0054368
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17=2.0664e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17=-2.0481e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17=0.0042182
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18=0.94584
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18=-0.0020089
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18=-0.0053067
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18=-0.0067852
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18=0.006337
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18=-8.4823e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18=-6.9974e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18=0.0031264
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19=0.65475
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19=-0.001468
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19=-0.0084439
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19=0.027564
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19=0.0050271
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19=-5.7219e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19=-3.4263e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19=0.24382
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20=0.40996
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20=-0.00057663
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20=-0.044961
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20=0.014184
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20=8.3656e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20=-1.5765e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20=-7260.8
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21=-4658.5
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21=0.2694
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21=-0.0022418
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21=-0.013905
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21=0.014513
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21=-2.0769e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21=-8.3428e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22=-0.026269
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22=-0.016505
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22=0.26022
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22=-0.0004019
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22=-0.039011
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22=-0.046788
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22=0.010589
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22=5.6891e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22=-3.7472e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23=0.00030057
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23=-0.00099596
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23=-0.030861
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23=0.0031886
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23=0.0055349
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23=1.0927e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23=-2.8385e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24=-7.2761e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24=0.0033354
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24=0.95716
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24=-0.0022322
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24=-0.010216
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24=-0.0055189
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24=0.0070116
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24=-3.9652e-13
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25=-3.0631e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25=-6.245e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25=0.0014436
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25=0.68151
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25=-0.0019888
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25=-0.011358
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25=0.0017263
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25=0.0051856
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26=0.01229
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26=8.1881e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26=-2.6025e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26=-4337.2
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26=-0.0012339
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26=-0.035371
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27=-0.030383
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27=0.014239
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27=4.5811e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27=-1.2254e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27=-2676.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27=0.21074
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27=-0.0035336
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28=0.19325
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28=-0.0026845
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28=-0.032078
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28=0.0103
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28=5.7493e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28=-9.5919e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28=-2381.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29=0.35973
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29=-0.0014642
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29=-0.018211
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29=-0.053694
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29=0.012737
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29=-3.3236e-15
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29=-4.07e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29=-0.030513
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30=0.072725
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30=-0.0010212
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30=-0.031
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30=0.0092162
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30=0.0059601
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30=3.7661e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30=-2.7739e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30=0.0059804
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31=0.92465
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31=-0.0022994
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31=-0.010998
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31=0.0025372
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31=0.0073413
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31=-1.9471e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31=-6.6952e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31=0.0015777
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32=0.65519
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32=-0.0019144
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32=-0.011028
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32=0.0024734
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32=0.0053534
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32=-2.3348e-14
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32=-5.6903e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32=0.0012195
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33=-4051.8
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33=0.5759
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33=-0.0018092
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33=-0.035798
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33=0.014803
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33=1.1162e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33=-5.3659e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34=-2166.3
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34=0.17738
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34=-0.0028276
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34=-0.024029
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34=0.010653
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34=1.1722e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34=-9.18e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35=-3.2583e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35=-0.0088062
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35=-1.9931e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35=5.2901e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35=0.33276
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35=-0.00038276
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35=-0.038399
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35=0.0034401
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35=-2.6122e-12
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36=-5.4782e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36=8.9661e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36=-1.729e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36=1.1815e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36=1.0031
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36=-0.00016769
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36=-0.020294
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36=0.0036381
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37=-0.00045955
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37=-2.7776e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37=1.4353e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37=-0.038852
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37=-1.0655e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37=6.8453e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37=0.29485
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37=0.00056132
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37=-0.019438
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38=-0.019654
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38=0.0022325
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38=8.4779e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38=2.9583e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38=-0.03654
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38=1.3015e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38=6.6762e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38=0.2561
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38=0.00070803
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39=0.57176
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39=-0.00024014
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39=-0.0060422
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39=0.0035435
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39=-6.323e-14
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39=1.287e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39=6.023e-9
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39=4.5041e-10
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40=0.19947
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40=-0.0033102
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40=0.026597
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40=0.012033
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40=-6.398e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40=-1.6127e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40=-8184.5
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41=0.00054213
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41=-0.040365
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41=0.0038952
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41=-2.8884e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41=-1.7185e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41=-2862.9
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42=0.29652
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42=-0.00074922
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42=-0.016885
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42=0.0080679
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42=7.3269e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42=-5.0772e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42=-758.34
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43=8.9949e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43=1.035e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43=0.19448
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43=-0.0016469
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43=-0.021918
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43=0.0088136
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43=-2.9651e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43=-8.0853e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44=6.6709e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44=3.901e-10
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44=0.31628
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44=-0.0021865
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44=-0.016043
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44=0.008385
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44=-2.8257e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44=-9.0212e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45=2.8576e-9
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45=3.2982e-11
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45=0.59252
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45=-0.00096288
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45=-0.01408
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45=0.0052573
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45=-3.9682e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45=-2.4517e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46=-9.1102e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46=-3564.6
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46=0.073602
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46=-0.0017827
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46=-0.0078965
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46=0.011489
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46=-3.6719e-12
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47=-1.0983e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47=-8.3074e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47=-3103.8
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47=0.19095
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47=-0.0024249
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47=-0.020135
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47=0.011567
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48=0.0074734
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48=-4.1147e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48=-7.9245e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48=-3508.2
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48=0.00035919
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48=-0.063256
.include "sky130_fd_pr__pfet_g5v0d10v5.pm3.spice"