* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param globalk=1
.param localkswitch=1
.param capunits='1.0*1e-6'
.param mcp1f_ca_w_0_150_s_0_210=1.06e-04
.param mcp1f_cc_w_0_150_s_0_210=7.62e-11
.param mcp1f_cf_w_0_150_s_0_210=1.03e-11
.param mcp1f_ca_w_0_150_s_0_263=1.06e-04
.param mcp1f_cc_w_0_150_s_0_263=6.19e-11
.param mcp1f_cf_w_0_150_s_0_263=1.25e-11
.param mcp1f_ca_w_0_150_s_0_315=1.06e-04
.param mcp1f_cc_w_0_150_s_0_315=5.27e-11
.param mcp1f_cf_w_0_150_s_0_315=1.45e-11
.param mcp1f_ca_w_0_150_s_0_420=1.06e-04
.param mcp1f_cc_w_0_150_s_0_420=4.04e-11
.param mcp1f_cf_w_0_150_s_0_420=1.85e-11
.param mcp1f_ca_w_0_150_s_0_525=1.06e-04
.param mcp1f_cc_w_0_150_s_0_525=3.29e-11
.param mcp1f_cf_w_0_150_s_0_525=2.17e-11
.param mcp1f_ca_w_0_150_s_0_630=1.06e-04
.param mcp1f_cc_w_0_150_s_0_630=2.76e-11
.param mcp1f_cf_w_0_150_s_0_630=2.46e-11
.param mcp1f_ca_w_0_150_s_0_840=1.06e-04
.param mcp1f_cc_w_0_150_s_0_840=2.03e-11
.param mcp1f_cf_w_0_150_s_0_840=2.94e-11
.param mcp1f_ca_w_0_150_s_1_260=1.06e-04
.param mcp1f_cc_w_0_150_s_1_260=1.18e-11
.param mcp1f_cf_w_0_150_s_1_260=3.62e-11
.param mcp1f_ca_w_0_150_s_2_310=1.06e-04
.param mcp1f_cc_w_0_150_s_2_310=5.10e-12
.param mcp1f_cf_w_0_150_s_2_310=4.24e-11
.param mcp1f_ca_w_0_150_s_5_250=1.06e-04
.param mcp1f_cc_w_0_150_s_5_250=1.20e-12
.param mcp1f_cf_w_0_150_s_5_250=4.63e-11
.param mcp1f_ca_w_1_200_s_0_210=1.06e-04
.param mcp1f_cc_w_1_200_s_0_210=9.44e-11
.param mcp1f_cf_w_1_200_s_0_210=1.02e-11
.param mcp1f_ca_w_1_200_s_0_263=1.06e-04
.param mcp1f_cc_w_1_200_s_0_263=7.89e-11
.param mcp1f_cf_w_1_200_s_0_263=1.25e-11
.param mcp1f_ca_w_1_200_s_0_315=1.06e-04
.param mcp1f_cc_w_1_200_s_0_315=6.86e-11
.param mcp1f_cf_w_1_200_s_0_315=1.46e-11
.param mcp1f_ca_w_1_200_s_0_420=1.06e-04
.param mcp1f_cc_w_1_200_s_0_420=5.49e-11
.param mcp1f_cf_w_1_200_s_0_420=1.84e-11
.param mcp1f_ca_w_1_200_s_0_525=1.06e-04
.param mcp1f_cc_w_1_200_s_0_525=4.61e-11
.param mcp1f_cf_w_1_200_s_0_525=2.19e-11
.param mcp1f_ca_w_1_200_s_0_630=1.06e-04
.param mcp1f_cc_w_1_200_s_0_630=3.98e-11
.param mcp1f_cf_w_1_200_s_0_630=2.49e-11
.param mcp1f_ca_w_1_200_s_0_840=1.06e-04
.param mcp1f_cc_w_1_200_s_0_840=3.12e-11
.param mcp1f_cf_w_1_200_s_0_840=2.99e-11
.param mcp1f_ca_w_1_200_s_1_260=1.06e-04
.param mcp1f_cc_w_1_200_s_1_260=2.14e-11
.param mcp1f_cf_w_1_200_s_1_260=3.71e-11
.param mcp1f_ca_w_1_200_s_2_310=1.06e-04
.param mcp1f_cc_w_1_200_s_2_310=1.08e-11
.param mcp1f_cf_w_1_200_s_2_310=4.64e-11
.param mcp1f_ca_w_1_200_s_5_250=1.06e-04
.param mcp1f_cc_w_1_200_s_5_250=3.40e-12
.param mcp1f_cf_w_1_200_s_5_250=5.36e-11
.param mcl1f_ca_w_0_170_s_0_180=3.69e-05
.param mcl1f_cc_w_0_170_s_0_180=7.98e-11
.param mcl1f_cf_w_0_170_s_0_180=3.26e-12
.param mcl1f_ca_w_0_170_s_0_225=3.69e-05
.param mcl1f_cc_w_0_170_s_0_225=6.83e-11
.param mcl1f_cf_w_0_170_s_0_225=4.04e-12
.param mcl1f_ca_w_0_170_s_0_270=3.69e-05
.param mcl1f_cc_w_0_170_s_0_270=6.07e-11
.param mcl1f_cf_w_0_170_s_0_270=4.81e-12
.param mcl1f_ca_w_0_170_s_0_360=3.69e-05
.param mcl1f_cc_w_0_170_s_0_360=4.97e-11
.param mcl1f_cf_w_0_170_s_0_360=6.42e-12
.param mcl1f_ca_w_0_170_s_0_450=3.69e-05
.param mcl1f_cc_w_0_170_s_0_450=4.29e-11
.param mcl1f_cf_w_0_170_s_0_450=7.78e-12
.param mcl1f_ca_w_0_170_s_0_540=3.69e-05
.param mcl1f_cc_w_0_170_s_0_540=3.73e-11
.param mcl1f_cf_w_0_170_s_0_540=9.40e-12
.param mcl1f_ca_w_0_170_s_0_720=3.69e-05
.param mcl1f_cc_w_0_170_s_0_720=3.01e-11
.param mcl1f_cf_w_0_170_s_0_720=1.20e-11
.param mcl1f_ca_w_0_170_s_1_080=3.69e-05
.param mcl1f_cc_w_0_170_s_1_080=2.13e-11
.param mcl1f_cf_w_0_170_s_1_080=1.66e-11
.param mcl1f_ca_w_0_170_s_1_980=3.69e-05
.param mcl1f_cc_w_0_170_s_1_980=1.14e-11
.param mcl1f_cf_w_0_170_s_1_980=2.36e-11
.param mcl1f_ca_w_0_170_s_4_500=3.69e-05
.param mcl1f_cc_w_0_170_s_4_500=3.41e-12
.param mcl1f_cf_w_0_170_s_4_500=3.09e-11
.param mcl1f_ca_w_1_360_s_0_180=3.69e-05
.param mcl1f_cc_w_1_360_s_0_180=1.02e-10
.param mcl1f_cf_w_1_360_s_0_180=3.26e-12
.param mcl1f_ca_w_1_360_s_0_225=3.69e-05
.param mcl1f_cc_w_1_360_s_0_225=8.88e-11
.param mcl1f_cf_w_1_360_s_0_225=4.04e-12
.param mcl1f_ca_w_1_360_s_0_270=3.69e-05
.param mcl1f_cc_w_1_360_s_0_270=7.95e-11
.param mcl1f_cf_w_1_360_s_0_270=4.82e-12
.param mcl1f_ca_w_1_360_s_0_360=3.69e-05
.param mcl1f_cc_w_1_360_s_0_360=6.68e-11
.param mcl1f_cf_w_1_360_s_0_360=6.35e-12
.param mcl1f_ca_w_1_360_s_0_450=3.69e-05
.param mcl1f_cc_w_1_360_s_0_450=5.83e-11
.param mcl1f_cf_w_1_360_s_0_450=7.83e-12
.param mcl1f_ca_w_1_360_s_0_540=3.69e-05
.param mcl1f_cc_w_1_360_s_0_540=5.20e-11
.param mcl1f_cf_w_1_360_s_0_540=9.25e-12
.param mcl1f_ca_w_1_360_s_0_720=3.69e-05
.param mcl1f_cc_w_1_360_s_0_720=4.31e-11
.param mcl1f_cf_w_1_360_s_0_720=1.19e-11
.param mcl1f_ca_w_1_360_s_1_080=3.69e-05
.param mcl1f_cc_w_1_360_s_1_080=3.23e-11
.param mcl1f_cf_w_1_360_s_1_080=1.67e-11
.param mcl1f_ca_w_1_360_s_1_980=3.69e-05
.param mcl1f_cc_w_1_360_s_1_980=1.90e-11
.param mcl1f_cf_w_1_360_s_1_980=2.53e-11
.param mcl1f_ca_w_1_360_s_4_500=3.69e-05
.param mcl1f_cc_w_1_360_s_4_500=7.05e-12
.param mcl1f_cf_w_1_360_s_4_500=3.57e-11
.param mcl1d_ca_w_0_170_s_0_180=5.53e-05
.param mcl1d_cc_w_0_170_s_0_180=7.74e-11
.param mcl1d_cf_w_0_170_s_0_180=4.83e-12
.param mcl1d_ca_w_0_170_s_0_225=5.53e-05
.param mcl1d_cc_w_0_170_s_0_225=6.56e-11
.param mcl1d_cf_w_0_170_s_0_225=5.98e-12
.param mcl1d_ca_w_0_170_s_0_270=5.53e-05
.param mcl1d_cc_w_0_170_s_0_270=5.78e-11
.param mcl1d_cf_w_0_170_s_0_270=7.08e-12
.param mcl1d_ca_w_0_170_s_0_360=5.53e-05
.param mcl1d_cc_w_0_170_s_0_360=4.66e-11
.param mcl1d_cf_w_0_170_s_0_360=9.37e-12
.param mcl1d_ca_w_0_170_s_0_450=5.53e-05
.param mcl1d_cc_w_0_170_s_0_450=3.96e-11
.param mcl1d_cf_w_0_170_s_0_450=1.13e-11
.param mcl1d_ca_w_0_170_s_0_540=5.53e-05
.param mcl1d_cc_w_0_170_s_0_540=3.39e-11
.param mcl1d_cf_w_0_170_s_0_540=1.35e-11
.param mcl1d_ca_w_0_170_s_0_720=5.53e-05
.param mcl1d_cc_w_0_170_s_0_720=2.64e-11
.param mcl1d_cf_w_0_170_s_0_720=1.70e-11
.param mcl1d_ca_w_0_170_s_1_080=5.53e-05
.param mcl1d_cc_w_0_170_s_1_080=1.75e-11
.param mcl1d_cf_w_0_170_s_1_080=2.25e-11
.param mcl1d_ca_w_0_170_s_1_980=5.53e-05
.param mcl1d_cc_w_0_170_s_1_980=8.42e-12
.param mcl1d_cf_w_0_170_s_1_980=3.00e-11
.param mcl1d_ca_w_0_170_s_4_500=5.53e-05
.param mcl1d_cc_w_0_170_s_4_500=2.28e-12
.param mcl1d_cf_w_0_170_s_4_500=3.59e-11
.param mcl1d_ca_w_1_360_s_0_180=5.53e-05
.param mcl1d_cc_w_1_360_s_0_180=9.72e-11
.param mcl1d_cf_w_1_360_s_0_180=4.83e-12
.param mcl1d_ca_w_1_360_s_0_225=5.53e-05
.param mcl1d_cc_w_1_360_s_0_225=8.44e-11
.param mcl1d_cf_w_1_360_s_0_225=5.98e-12
.param mcl1d_ca_w_1_360_s_0_270=5.53e-05
.param mcl1d_cc_w_1_360_s_0_270=7.51e-11
.param mcl1d_cf_w_1_360_s_0_270=7.11e-12
.param mcl1d_ca_w_1_360_s_0_360=5.53e-05
.param mcl1d_cc_w_1_360_s_0_360=6.24e-11
.param mcl1d_cf_w_1_360_s_0_360=9.29e-12
.param mcl1d_ca_w_1_360_s_0_450=5.53e-05
.param mcl1d_cc_w_1_360_s_0_450=5.39e-11
.param mcl1d_cf_w_1_360_s_0_450=1.14e-11
.param mcl1d_ca_w_1_360_s_0_540=5.53e-05
.param mcl1d_cc_w_1_360_s_0_540=4.76e-11
.param mcl1d_cf_w_1_360_s_0_540=1.33e-11
.param mcl1d_ca_w_1_360_s_0_720=5.53e-05
.param mcl1d_cc_w_1_360_s_0_720=3.87e-11
.param mcl1d_cf_w_1_360_s_0_720=1.70e-11
.param mcl1d_ca_w_1_360_s_1_080=5.53e-05
.param mcl1d_cc_w_1_360_s_1_080=2.80e-11
.param mcl1d_cf_w_1_360_s_1_080=2.29e-11
.param mcl1d_ca_w_1_360_s_1_980=5.53e-05
.param mcl1d_cc_w_1_360_s_1_980=1.55e-11
.param mcl1d_cf_w_1_360_s_1_980=3.25e-11
.param mcl1d_ca_w_1_360_s_4_500=5.53e-05
.param mcl1d_cc_w_1_360_s_4_500=5.35e-12
.param mcl1d_cf_w_1_360_s_4_500=4.19e-11
.param mcl1p1_ca_w_0_170_s_0_180=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_180=7.32e-11
.param mcl1p1_cf_w_0_170_s_0_180=8.06e-12
.param mcl1p1_ca_w_0_170_s_0_225=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_225=6.12e-11
.param mcl1p1_cf_w_0_170_s_0_225=9.91e-12
.param mcl1p1_ca_w_0_170_s_0_270=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_270=5.32e-11
.param mcl1p1_cf_w_0_170_s_0_270=1.17e-11
.param mcl1p1_ca_w_0_170_s_0_360=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_360=4.16e-11
.param mcl1p1_cf_w_0_170_s_0_360=1.52e-11
.param mcl1p1_ca_w_0_170_s_0_450=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_450=3.45e-11
.param mcl1p1_cf_w_0_170_s_0_450=1.80e-11
.param mcl1p1_ca_w_0_170_s_0_540=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_540=2.86e-11
.param mcl1p1_cf_w_0_170_s_0_540=2.12e-11
.param mcl1p1_ca_w_0_170_s_0_720=9.41e-05
.param mcl1p1_cc_w_0_170_s_0_720=2.11e-11
.param mcl1p1_cf_w_0_170_s_0_720=2.58e-11
.param mcl1p1_ca_w_0_170_s_1_080=9.41e-05
.param mcl1p1_cc_w_0_170_s_1_080=1.28e-11
.param mcl1p1_cf_w_0_170_s_1_080=3.22e-11
.param mcl1p1_ca_w_0_170_s_1_980=9.41e-05
.param mcl1p1_cc_w_0_170_s_1_980=5.43e-12
.param mcl1p1_cf_w_0_170_s_1_980=3.89e-11
.param mcl1p1_ca_w_0_170_s_4_500=9.41e-05
.param mcl1p1_cc_w_0_170_s_4_500=1.35e-12
.param mcl1p1_cf_w_0_170_s_4_500=4.29e-11
.param mcl1p1_ca_w_1_360_s_0_180=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_180=9.13e-11
.param mcl1p1_cf_w_1_360_s_0_180=8.11e-12
.param mcl1p1_ca_w_1_360_s_0_225=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_225=7.85e-11
.param mcl1p1_cf_w_1_360_s_0_225=9.97e-12
.param mcl1p1_ca_w_1_360_s_0_270=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_270=6.93e-11
.param mcl1p1_cf_w_1_360_s_0_270=1.18e-11
.param mcl1p1_ca_w_1_360_s_0_360=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_360=5.66e-11
.param mcl1p1_cf_w_1_360_s_0_360=1.51e-11
.param mcl1p1_ca_w_1_360_s_0_450=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_450=4.82e-11
.param mcl1p1_cf_w_1_360_s_0_450=1.82e-11
.param mcl1p1_ca_w_1_360_s_0_540=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_540=4.19e-11
.param mcl1p1_cf_w_1_360_s_0_540=2.11e-11
.param mcl1p1_ca_w_1_360_s_0_720=9.41e-05
.param mcl1p1_cc_w_1_360_s_0_720=3.32e-11
.param mcl1p1_cf_w_1_360_s_0_720=2.59e-11
.param mcl1p1_ca_w_1_360_s_1_080=9.41e-05
.param mcl1p1_cc_w_1_360_s_1_080=2.31e-11
.param mcl1p1_cf_w_1_360_s_1_080=3.31e-11
.param mcl1p1_ca_w_1_360_s_1_980=9.41e-05
.param mcl1p1_cc_w_1_360_s_1_980=1.19e-11
.param mcl1p1_cf_w_1_360_s_1_980=4.28e-11
.param mcl1p1_ca_w_1_360_s_4_500=9.41e-05
.param mcl1p1_cc_w_1_360_s_4_500=3.90e-12
.param mcl1p1_cf_w_1_360_s_4_500=5.06e-11
.param mcm1f_ca_w_0_140_s_0_140=2.58e-05
.param mcm1f_cc_w_0_140_s_0_140=1.05e-10
.param mcm1f_cf_w_0_140_s_0_140=1.79e-12
.param mcm1f_ca_w_0_140_s_0_175=2.58e-05
.param mcm1f_cc_w_0_140_s_0_175=1.03e-10
.param mcm1f_cf_w_0_140_s_0_175=2.23e-12
.param mcm1f_ca_w_0_140_s_0_210=2.58e-05
.param mcm1f_cc_w_0_140_s_0_210=9.77e-11
.param mcm1f_cf_w_0_140_s_0_210=2.68e-12
.param mcm1f_ca_w_0_140_s_0_280=2.58e-05
.param mcm1f_cc_w_0_140_s_0_280=8.76e-11
.param mcm1f_cf_w_0_140_s_0_280=3.56e-12
.param mcm1f_ca_w_0_140_s_0_350=2.58e-05
.param mcm1f_cc_w_0_140_s_0_350=7.63e-11
.param mcm1f_cf_w_0_140_s_0_350=4.42e-12
.param mcm1f_ca_w_0_140_s_0_420=2.58e-05
.param mcm1f_cc_w_0_140_s_0_420=6.70e-11
.param mcm1f_cf_w_0_140_s_0_420=5.31e-12
.param mcm1f_ca_w_0_140_s_0_560=2.58e-05
.param mcm1f_cc_w_0_140_s_0_560=5.45e-11
.param mcm1f_cf_w_0_140_s_0_560=6.93e-12
.param mcm1f_ca_w_0_140_s_0_840=2.58e-05
.param mcm1f_cc_w_0_140_s_0_840=4.05e-11
.param mcm1f_cf_w_0_140_s_0_840=1.00e-11
.param mcm1f_ca_w_0_140_s_1_540=2.58e-05
.param mcm1f_cc_w_0_140_s_1_540=2.47e-11
.param mcm1f_cf_w_0_140_s_1_540=1.65e-11
.param mcm1f_ca_w_0_140_s_3_500=2.58e-05
.param mcm1f_cc_w_0_140_s_3_500=1.00e-11
.param mcm1f_cf_w_0_140_s_3_500=2.70e-11
.param mcm1f_ca_w_1_120_s_0_140=2.58e-05
.param mcm1f_cc_w_1_120_s_0_140=1.31e-10
.param mcm1f_cf_w_1_120_s_0_140=1.82e-12
.param mcm1f_ca_w_1_120_s_0_175=2.58e-05
.param mcm1f_cc_w_1_120_s_0_175=1.27e-10
.param mcm1f_cf_w_1_120_s_0_175=2.28e-12
.param mcm1f_ca_w_1_120_s_0_210=2.58e-05
.param mcm1f_cc_w_1_120_s_0_210=1.21e-10
.param mcm1f_cf_w_1_120_s_0_210=2.72e-12
.param mcm1f_ca_w_1_120_s_0_280=2.58e-05
.param mcm1f_cc_w_1_120_s_0_280=1.07e-10
.param mcm1f_cf_w_1_120_s_0_280=3.61e-12
.param mcm1f_ca_w_1_120_s_0_350=2.58e-05
.param mcm1f_cc_w_1_120_s_0_350=9.46e-11
.param mcm1f_cf_w_1_120_s_0_350=4.47e-12
.param mcm1f_ca_w_1_120_s_0_420=2.58e-05
.param mcm1f_cc_w_1_120_s_0_420=8.38e-11
.param mcm1f_cf_w_1_120_s_0_420=5.33e-12
.param mcm1f_ca_w_1_120_s_0_560=2.58e-05
.param mcm1f_cc_w_1_120_s_0_560=6.88e-11
.param mcm1f_cf_w_1_120_s_0_560=6.98e-12
.param mcm1f_ca_w_1_120_s_0_840=2.58e-05
.param mcm1f_cc_w_1_120_s_0_840=5.20e-11
.param mcm1f_cf_w_1_120_s_0_840=1.01e-11
.param mcm1f_ca_w_1_120_s_1_540=2.58e-05
.param mcm1f_cc_w_1_120_s_1_540=3.29e-11
.param mcm1f_cf_w_1_120_s_1_540=1.69e-11
.param mcm1f_ca_w_1_120_s_3_500=2.58e-05
.param mcm1f_cc_w_1_120_s_3_500=1.47e-11
.param mcm1f_cf_w_1_120_s_3_500=2.88e-11
.param mcm1d_ca_w_0_140_s_0_140=3.36e-05
.param mcm1d_cc_w_0_140_s_0_140=1.04e-10
.param mcm1d_cf_w_0_140_s_0_140=2.32e-12
.param mcm1d_ca_w_0_140_s_0_175=3.36e-05
.param mcm1d_cc_w_0_140_s_0_175=1.02e-10
.param mcm1d_cf_w_0_140_s_0_175=2.90e-12
.param mcm1d_ca_w_0_140_s_0_210=3.36e-05
.param mcm1d_cc_w_0_140_s_0_210=9.66e-11
.param mcm1d_cf_w_0_140_s_0_210=3.49e-12
.param mcm1d_ca_w_0_140_s_0_280=3.36e-05
.param mcm1d_cc_w_0_140_s_0_280=8.60e-11
.param mcm1d_cf_w_0_140_s_0_280=4.62e-12
.param mcm1d_ca_w_0_140_s_0_350=3.36e-05
.param mcm1d_cc_w_0_140_s_0_350=7.46e-11
.param mcm1d_cf_w_0_140_s_0_350=5.73e-12
.param mcm1d_ca_w_0_140_s_0_420=3.36e-05
.param mcm1d_cc_w_0_140_s_0_420=6.53e-11
.param mcm1d_cf_w_0_140_s_0_420=6.87e-12
.param mcm1d_ca_w_0_140_s_0_560=3.36e-05
.param mcm1d_cc_w_0_140_s_0_560=5.27e-11
.param mcm1d_cf_w_0_140_s_0_560=8.91e-12
.param mcm1d_ca_w_0_140_s_0_840=3.36e-05
.param mcm1d_cc_w_0_140_s_0_840=3.84e-11
.param mcm1d_cf_w_0_140_s_0_840=1.28e-11
.param mcm1d_ca_w_0_140_s_1_540=3.36e-05
.param mcm1d_cc_w_0_140_s_1_540=2.23e-11
.param mcm1d_cf_w_0_140_s_1_540=2.05e-11
.param mcm1d_ca_w_0_140_s_3_500=3.36e-05
.param mcm1d_cc_w_0_140_s_3_500=8.26e-12
.param mcm1d_cf_w_0_140_s_3_500=3.15e-11
.param mcm1d_ca_w_1_120_s_0_140=3.36e-05
.param mcm1d_cc_w_1_120_s_0_140=1.28e-10
.param mcm1d_cf_w_1_120_s_0_140=2.39e-12
.param mcm1d_ca_w_1_120_s_0_175=3.36e-05
.param mcm1d_cc_w_1_120_s_0_175=1.24e-10
.param mcm1d_cf_w_1_120_s_0_175=2.96e-12
.param mcm1d_ca_w_1_120_s_0_210=3.36e-05
.param mcm1d_cc_w_1_120_s_0_210=1.18e-10
.param mcm1d_cf_w_1_120_s_0_210=3.54e-12
.param mcm1d_ca_w_1_120_s_0_280=3.36e-05
.param mcm1d_cc_w_1_120_s_0_280=1.04e-10
.param mcm1d_cf_w_1_120_s_0_280=4.68e-12
.param mcm1d_ca_w_1_120_s_0_350=3.36e-05
.param mcm1d_cc_w_1_120_s_0_350=9.17e-11
.param mcm1d_cf_w_1_120_s_0_350=5.80e-12
.param mcm1d_ca_w_1_120_s_0_420=3.36e-05
.param mcm1d_cc_w_1_120_s_0_420=8.11e-11
.param mcm1d_cf_w_1_120_s_0_420=6.89e-12
.param mcm1d_ca_w_1_120_s_0_560=3.36e-05
.param mcm1d_cc_w_1_120_s_0_560=6.60e-11
.param mcm1d_cf_w_1_120_s_0_560=8.99e-12
.param mcm1d_ca_w_1_120_s_0_840=3.36e-05
.param mcm1d_cc_w_1_120_s_0_840=4.91e-11
.param mcm1d_cf_w_1_120_s_0_840=1.29e-11
.param mcm1d_ca_w_1_120_s_1_540=3.36e-05
.param mcm1d_cc_w_1_120_s_1_540=3.01e-11
.param mcm1d_cf_w_1_120_s_1_540=2.09e-11
.param mcm1d_ca_w_1_120_s_3_500=3.36e-05
.param mcm1d_cc_w_1_120_s_3_500=1.26e-11
.param mcm1d_cf_w_1_120_s_3_500=3.36e-11
.param mcm1p1_ca_w_0_140_s_0_140=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_140=1.03e-10
.param mcm1p1_cf_w_0_140_s_0_140=3.09e-12
.param mcm1p1_ca_w_0_140_s_0_175=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_175=1.01e-10
.param mcm1p1_cf_w_0_140_s_0_175=3.87e-12
.param mcm1p1_ca_w_0_140_s_0_210=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_210=9.50e-11
.param mcm1p1_cf_w_0_140_s_0_210=4.64e-12
.param mcm1p1_ca_w_0_140_s_0_280=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_280=8.43e-11
.param mcm1p1_cf_w_0_140_s_0_280=6.14e-12
.param mcm1p1_ca_w_0_140_s_0_350=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_350=7.26e-11
.param mcm1p1_cf_w_0_140_s_0_350=7.60e-12
.param mcm1p1_ca_w_0_140_s_0_420=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_420=6.31e-11
.param mcm1p1_cf_w_0_140_s_0_420=9.06e-12
.param mcm1p1_ca_w_0_140_s_0_560=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_560=5.03e-11
.param mcm1p1_cf_w_0_140_s_0_560=1.17e-11
.param mcm1p1_ca_w_0_140_s_0_840=4.48e-05
.param mcm1p1_cc_w_0_140_s_0_840=3.57e-11
.param mcm1p1_cf_w_0_140_s_0_840=1.65e-11
.param mcm1p1_ca_w_0_140_s_1_540=4.48e-05
.param mcm1p1_cc_w_0_140_s_1_540=1.96e-11
.param mcm1p1_cf_w_0_140_s_1_540=2.55e-11
.param mcm1p1_ca_w_0_140_s_3_500=4.48e-05
.param mcm1p1_cc_w_0_140_s_3_500=6.59e-12
.param mcm1p1_cf_w_0_140_s_3_500=3.65e-11
.param mcm1p1_ca_w_1_120_s_0_140=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_140=1.25e-10
.param mcm1p1_cf_w_1_120_s_0_140=3.22e-12
.param mcm1p1_ca_w_1_120_s_0_175=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_175=1.21e-10
.param mcm1p1_cf_w_1_120_s_0_175=4.00e-12
.param mcm1p1_ca_w_1_120_s_0_210=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_210=1.14e-10
.param mcm1p1_cf_w_1_120_s_0_210=4.77e-12
.param mcm1p1_ca_w_1_120_s_0_280=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_280=1.01e-10
.param mcm1p1_cf_w_1_120_s_0_280=6.26e-12
.param mcm1p1_ca_w_1_120_s_0_350=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_350=8.83e-11
.param mcm1p1_cf_w_1_120_s_0_350=7.72e-12
.param mcm1p1_ca_w_1_120_s_0_420=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_420=7.77e-11
.param mcm1p1_cf_w_1_120_s_0_420=9.16e-12
.param mcm1p1_ca_w_1_120_s_0_560=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_560=6.27e-11
.param mcm1p1_cf_w_1_120_s_0_560=1.18e-11
.param mcm1p1_ca_w_1_120_s_0_840=4.48e-05
.param mcm1p1_cc_w_1_120_s_0_840=4.59e-11
.param mcm1p1_cf_w_1_120_s_0_840=1.68e-11
.param mcm1p1_ca_w_1_120_s_1_540=4.48e-05
.param mcm1p1_cc_w_1_120_s_1_540=2.71e-11
.param mcm1p1_cf_w_1_120_s_1_540=2.61e-11
.param mcm1p1_ca_w_1_120_s_3_500=4.48e-05
.param mcm1p1_cc_w_1_120_s_3_500=1.07e-11
.param mcm1p1_cf_w_1_120_s_3_500=3.92e-11
.param mcm1l1_ca_w_0_140_s_0_140=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_140=9.58e-11
.param mcm1l1_cf_w_0_140_s_0_140=7.43e-12
.param mcm1l1_ca_w_0_140_s_0_175=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_175=9.38e-11
.param mcm1l1_cf_w_0_140_s_0_175=9.39e-12
.param mcm1l1_ca_w_0_140_s_0_210=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_210=8.80e-11
.param mcm1l1_cf_w_0_140_s_0_210=1.13e-11
.param mcm1l1_ca_w_0_140_s_0_280=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_280=7.59e-11
.param mcm1l1_cf_w_0_140_s_0_280=1.48e-11
.param mcm1l1_ca_w_0_140_s_0_350=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_350=6.44e-11
.param mcm1l1_cf_w_0_140_s_0_350=1.81e-11
.param mcm1l1_ca_w_0_140_s_0_420=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_420=5.44e-11
.param mcm1l1_cf_w_0_140_s_0_420=2.12e-11
.param mcm1l1_ca_w_0_140_s_0_560=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_560=4.13e-11
.param mcm1l1_cf_w_0_140_s_0_560=2.65e-11
.param mcm1l1_ca_w_0_140_s_0_840=1.14e-04
.param mcm1l1_cc_w_0_140_s_0_840=2.70e-11
.param mcm1l1_cf_w_0_140_s_0_840=3.47e-11
.param mcm1l1_ca_w_0_140_s_1_540=1.14e-04
.param mcm1l1_cc_w_0_140_s_1_540=1.25e-11
.param mcm1l1_cf_w_0_140_s_1_540=4.62e-11
.param mcm1l1_ca_w_0_140_s_3_500=1.14e-04
.param mcm1l1_cc_w_0_140_s_3_500=3.55e-12
.param mcm1l1_cf_w_0_140_s_3_500=5.51e-11
.param mcm1l1_ca_w_1_120_s_0_140=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_140=1.15e-10
.param mcm1l1_cf_w_1_120_s_0_140=7.56e-12
.param mcm1l1_ca_w_1_120_s_0_175=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_175=1.10e-10
.param mcm1l1_cf_w_1_120_s_0_175=9.50e-12
.param mcm1l1_ca_w_1_120_s_0_210=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_210=1.04e-10
.param mcm1l1_cf_w_1_120_s_0_210=1.14e-11
.param mcm1l1_ca_w_1_120_s_0_280=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_280=9.04e-11
.param mcm1l1_cf_w_1_120_s_0_280=1.49e-11
.param mcm1l1_ca_w_1_120_s_0_350=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_350=7.72e-11
.param mcm1l1_cf_w_1_120_s_0_350=1.82e-11
.param mcm1l1_ca_w_1_120_s_0_420=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_420=6.73e-11
.param mcm1l1_cf_w_1_120_s_0_420=2.13e-11
.param mcm1l1_ca_w_1_120_s_0_560=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_560=5.26e-11
.param mcm1l1_cf_w_1_120_s_0_560=2.66e-11
.param mcm1l1_ca_w_1_120_s_0_840=1.14e-04
.param mcm1l1_cc_w_1_120_s_0_840=3.64e-11
.param mcm1l1_cf_w_1_120_s_0_840=3.50e-11
.param mcm1l1_ca_w_1_120_s_1_540=1.14e-04
.param mcm1l1_cc_w_1_120_s_1_540=1.97e-11
.param mcm1l1_cf_w_1_120_s_1_540=4.74e-11
.param mcm1l1_ca_w_1_120_s_3_500=1.14e-04
.param mcm1l1_cc_w_1_120_s_3_500=7.00e-12
.param mcm1l1_cf_w_1_120_s_3_500=5.94e-11
.param mcm2f_ca_w_0_140_s_0_140=1.75e-05
.param mcm2f_cc_w_0_140_s_0_140=1.07e-10
.param mcm2f_cf_w_0_140_s_0_140=1.22e-12
.param mcm2f_ca_w_0_140_s_0_175=1.75e-05
.param mcm2f_cc_w_0_140_s_0_175=1.04e-10
.param mcm2f_cf_w_0_140_s_0_175=1.53e-12
.param mcm2f_ca_w_0_140_s_0_210=1.75e-05
.param mcm2f_cc_w_0_140_s_0_210=9.87e-11
.param mcm2f_cf_w_0_140_s_0_210=1.84e-12
.param mcm2f_ca_w_0_140_s_0_280=1.75e-05
.param mcm2f_cc_w_0_140_s_0_280=8.88e-11
.param mcm2f_cf_w_0_140_s_0_280=2.44e-12
.param mcm2f_ca_w_0_140_s_0_350=1.75e-05
.param mcm2f_cc_w_0_140_s_0_350=7.76e-11
.param mcm2f_cf_w_0_140_s_0_350=3.03e-12
.param mcm2f_ca_w_0_140_s_0_420=1.75e-05
.param mcm2f_cc_w_0_140_s_0_420=6.85e-11
.param mcm2f_cf_w_0_140_s_0_420=3.65e-12
.param mcm2f_ca_w_0_140_s_0_560=1.75e-05
.param mcm2f_cc_w_0_140_s_0_560=5.62e-11
.param mcm2f_cf_w_0_140_s_0_560=4.77e-12
.param mcm2f_ca_w_0_140_s_0_840=1.75e-05
.param mcm2f_cc_w_0_140_s_0_840=4.26e-11
.param mcm2f_cf_w_0_140_s_0_840=6.98e-12
.param mcm2f_ca_w_0_140_s_1_540=1.75e-05
.param mcm2f_cc_w_0_140_s_1_540=2.74e-11
.param mcm2f_cf_w_0_140_s_1_540=1.19e-11
.param mcm2f_ca_w_0_140_s_3_500=1.75e-05
.param mcm2f_cc_w_0_140_s_3_500=1.27e-11
.param mcm2f_cf_w_0_140_s_3_500=2.10e-11
.param mcm2f_ca_w_1_120_s_0_140=1.75e-05
.param mcm2f_cc_w_1_120_s_0_140=1.33e-10
.param mcm2f_cf_w_1_120_s_0_140=1.25e-12
.param mcm2f_ca_w_1_120_s_0_175=1.75e-05
.param mcm2f_cc_w_1_120_s_0_175=1.29e-10
.param mcm2f_cf_w_1_120_s_0_175=1.55e-12
.param mcm2f_ca_w_1_120_s_0_210=1.75e-05
.param mcm2f_cc_w_1_120_s_0_210=1.23e-10
.param mcm2f_cf_w_1_120_s_0_210=1.86e-12
.param mcm2f_ca_w_1_120_s_0_280=1.75e-05
.param mcm2f_cc_w_1_120_s_0_280=1.10e-10
.param mcm2f_cf_w_1_120_s_0_280=2.47e-12
.param mcm2f_ca_w_1_120_s_0_350=1.75e-05
.param mcm2f_cc_w_1_120_s_0_350=9.70e-11
.param mcm2f_cf_w_1_120_s_0_350=3.06e-12
.param mcm2f_ca_w_1_120_s_0_420=1.75e-05
.param mcm2f_cc_w_1_120_s_0_420=8.65e-11
.param mcm2f_cf_w_1_120_s_0_420=3.66e-12
.param mcm2f_ca_w_1_120_s_0_560=1.75e-05
.param mcm2f_cc_w_1_120_s_0_560=7.16e-11
.param mcm2f_cf_w_1_120_s_0_560=4.81e-12
.param mcm2f_ca_w_1_120_s_0_840=1.75e-05
.param mcm2f_cc_w_1_120_s_0_840=5.50e-11
.param mcm2f_cf_w_1_120_s_0_840=7.06e-12
.param mcm2f_ca_w_1_120_s_1_540=1.75e-05
.param mcm2f_cc_w_1_120_s_1_540=3.62e-11
.param mcm2f_cf_w_1_120_s_1_540=1.21e-11
.param mcm2f_ca_w_1_120_s_3_500=1.75e-05
.param mcm2f_cc_w_1_120_s_3_500=1.79e-11
.param mcm2f_cf_w_1_120_s_3_500=2.22e-11
.param mcm2d_ca_w_0_140_s_0_140=2.08e-05
.param mcm2d_cc_w_0_140_s_0_140=1.05e-10
.param mcm2d_cf_w_0_140_s_0_140=1.45e-12
.param mcm2d_ca_w_0_140_s_0_175=2.08e-05
.param mcm2d_cc_w_0_140_s_0_175=1.03e-10
.param mcm2d_cf_w_0_140_s_0_175=1.81e-12
.param mcm2d_ca_w_0_140_s_0_210=2.08e-05
.param mcm2d_cc_w_0_140_s_0_210=9.82e-11
.param mcm2d_cf_w_0_140_s_0_210=2.18e-12
.param mcm2d_ca_w_0_140_s_0_280=2.08e-05
.param mcm2d_cc_w_0_140_s_0_280=8.83e-11
.param mcm2d_cf_w_0_140_s_0_280=2.89e-12
.param mcm2d_ca_w_0_140_s_0_350=2.08e-05
.param mcm2d_cc_w_0_140_s_0_350=7.70e-11
.param mcm2d_cf_w_0_140_s_0_350=3.59e-12
.param mcm2d_ca_w_0_140_s_0_420=2.08e-05
.param mcm2d_cc_w_0_140_s_0_420=6.74e-11
.param mcm2d_cf_w_0_140_s_0_420=4.32e-12
.param mcm2d_ca_w_0_140_s_0_560=2.08e-05
.param mcm2d_cc_w_0_140_s_0_560=5.52e-11
.param mcm2d_cf_w_0_140_s_0_560=5.62e-12
.param mcm2d_ca_w_0_140_s_0_840=2.08e-05
.param mcm2d_cc_w_0_140_s_0_840=4.16e-11
.param mcm2d_cf_w_0_140_s_0_840=8.21e-12
.param mcm2d_ca_w_0_140_s_1_540=2.08e-05
.param mcm2d_cc_w_0_140_s_1_540=2.60e-11
.param mcm2d_cf_w_0_140_s_1_540=1.37e-11
.param mcm2d_ca_w_0_140_s_3_500=2.08e-05
.param mcm2d_cc_w_0_140_s_3_500=1.14e-11
.param mcm2d_cf_w_0_140_s_3_500=2.35e-11
.param mcm2d_ca_w_1_120_s_0_140=2.08e-05
.param mcm2d_cc_w_1_120_s_0_140=1.32e-10
.param mcm2d_cf_w_1_120_s_0_140=1.49e-12
.param mcm2d_ca_w_1_120_s_0_175=2.08e-05
.param mcm2d_cc_w_1_120_s_0_175=1.28e-10
.param mcm2d_cf_w_1_120_s_0_175=1.85e-12
.param mcm2d_ca_w_1_120_s_0_210=2.08e-05
.param mcm2d_cc_w_1_120_s_0_210=1.22e-10
.param mcm2d_cf_w_1_120_s_0_210=2.21e-12
.param mcm2d_ca_w_1_120_s_0_280=2.08e-05
.param mcm2d_cc_w_1_120_s_0_280=1.08e-10
.param mcm2d_cf_w_1_120_s_0_280=2.92e-12
.param mcm2d_ca_w_1_120_s_0_350=2.08e-05
.param mcm2d_cc_w_1_120_s_0_350=9.54e-11
.param mcm2d_cf_w_1_120_s_0_350=3.63e-12
.param mcm2d_ca_w_1_120_s_0_420=2.08e-05
.param mcm2d_cc_w_1_120_s_0_420=8.50e-11
.param mcm2d_cf_w_1_120_s_0_420=4.32e-12
.param mcm2d_ca_w_1_120_s_0_560=2.08e-05
.param mcm2d_cc_w_1_120_s_0_560=7.00e-11
.param mcm2d_cf_w_1_120_s_0_560=5.68e-12
.param mcm2d_ca_w_1_120_s_0_840=2.08e-05
.param mcm2d_cc_w_1_120_s_0_840=5.33e-11
.param mcm2d_cf_w_1_120_s_0_840=8.27e-12
.param mcm2d_ca_w_1_120_s_1_540=2.08e-05
.param mcm2d_cc_w_1_120_s_1_540=3.45e-11
.param mcm2d_cf_w_1_120_s_1_540=1.40e-11
.param mcm2d_ca_w_1_120_s_3_500=2.08e-05
.param mcm2d_cc_w_1_120_s_3_500=1.63e-11
.param mcm2d_cf_w_1_120_s_3_500=2.50e-11
.param mcm2p1_ca_w_0_140_s_0_140=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_140=1.05e-10
.param mcm2p1_cf_w_0_140_s_0_140=1.72e-12
.param mcm2p1_ca_w_0_140_s_0_175=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_175=1.03e-10
.param mcm2p1_cf_w_0_140_s_0_175=2.14e-12
.param mcm2p1_ca_w_0_140_s_0_210=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_210=9.77e-11
.param mcm2p1_cf_w_0_140_s_0_210=2.58e-12
.param mcm2p1_ca_w_0_140_s_0_280=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_280=8.77e-11
.param mcm2p1_cf_w_0_140_s_0_280=3.42e-12
.param mcm2p1_ca_w_0_140_s_0_350=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_350=7.60e-11
.param mcm2p1_cf_w_0_140_s_0_350=4.24e-12
.param mcm2p1_ca_w_0_140_s_0_420=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_420=6.66e-11
.param mcm2p1_cf_w_0_140_s_0_420=5.10e-12
.param mcm2p1_ca_w_0_140_s_0_560=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_560=5.44e-11
.param mcm2p1_cf_w_0_140_s_0_560=6.65e-12
.param mcm2p1_ca_w_0_140_s_0_840=2.47e-05
.param mcm2p1_cc_w_0_140_s_0_840=4.04e-11
.param mcm2p1_cf_w_0_140_s_0_840=9.62e-12
.param mcm2p1_ca_w_0_140_s_1_540=2.47e-05
.param mcm2p1_cc_w_0_140_s_1_540=2.46e-11
.param mcm2p1_cf_w_0_140_s_1_540=1.59e-11
.param mcm2p1_ca_w_0_140_s_3_500=2.47e-05
.param mcm2p1_cc_w_0_140_s_3_500=1.01e-11
.param mcm2p1_cf_w_0_140_s_3_500=2.62e-11
.param mcm2p1_ca_w_1_120_s_0_140=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_140=1.30e-10
.param mcm2p1_cf_w_1_120_s_0_140=1.78e-12
.param mcm2p1_ca_w_1_120_s_0_175=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_175=1.26e-10
.param mcm2p1_cf_w_1_120_s_0_175=2.21e-12
.param mcm2p1_ca_w_1_120_s_0_210=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_210=1.20e-10
.param mcm2p1_cf_w_1_120_s_0_210=2.64e-12
.param mcm2p1_ca_w_1_120_s_0_280=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_280=1.07e-10
.param mcm2p1_cf_w_1_120_s_0_280=3.48e-12
.param mcm2p1_ca_w_1_120_s_0_350=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_350=9.38e-11
.param mcm2p1_cf_w_1_120_s_0_350=4.31e-12
.param mcm2p1_ca_w_1_120_s_0_420=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_420=8.32e-11
.param mcm2p1_cf_w_1_120_s_0_420=5.14e-12
.param mcm2p1_ca_w_1_120_s_0_560=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_560=6.85e-11
.param mcm2p1_cf_w_1_120_s_0_560=6.72e-12
.param mcm2p1_ca_w_1_120_s_0_840=2.47e-05
.param mcm2p1_cc_w_1_120_s_0_840=5.16e-11
.param mcm2p1_cf_w_1_120_s_0_840=9.73e-12
.param mcm2p1_ca_w_1_120_s_1_540=2.47e-05
.param mcm2p1_cc_w_1_120_s_1_540=3.27e-11
.param mcm2p1_cf_w_1_120_s_1_540=1.62e-11
.param mcm2p1_ca_w_1_120_s_3_500=2.47e-05
.param mcm2p1_cc_w_1_120_s_3_500=1.48e-11
.param mcm2p1_cf_w_1_120_s_3_500=2.79e-11
.param mcm2l1_ca_w_0_140_s_0_140=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_140=1.03e-10
.param mcm2l1_cf_w_0_140_s_0_140=2.54e-12
.param mcm2l1_ca_w_0_140_s_0_175=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_175=1.02e-10
.param mcm2l1_cf_w_0_140_s_0_175=3.18e-12
.param mcm2l1_ca_w_0_140_s_0_210=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_210=9.62e-11
.param mcm2l1_cf_w_0_140_s_0_210=3.83e-12
.param mcm2l1_ca_w_0_140_s_0_280=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_280=8.51e-11
.param mcm2l1_cf_w_0_140_s_0_280=5.07e-12
.param mcm2l1_ca_w_0_140_s_0_350=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_350=7.38e-11
.param mcm2l1_cf_w_0_140_s_0_350=6.28e-12
.param mcm2l1_ca_w_0_140_s_0_420=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_420=6.44e-11
.param mcm2l1_cf_w_0_140_s_0_420=7.51e-12
.param mcm2l1_ca_w_0_140_s_0_560=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_560=5.15e-11
.param mcm2l1_cf_w_0_140_s_0_560=9.75e-12
.param mcm2l1_ca_w_0_140_s_0_840=3.70e-05
.param mcm2l1_cc_w_0_140_s_0_840=3.71e-11
.param mcm2l1_cf_w_0_140_s_0_840=1.38e-11
.param mcm2l1_ca_w_0_140_s_1_540=3.70e-05
.param mcm2l1_cc_w_0_140_s_1_540=2.11e-11
.param mcm2l1_cf_w_0_140_s_1_540=2.20e-11
.param mcm2l1_ca_w_0_140_s_3_500=3.70e-05
.param mcm2l1_cc_w_0_140_s_3_500=7.54e-12
.param mcm2l1_cf_w_0_140_s_3_500=3.29e-11
.param mcm2l1_ca_w_1_120_s_0_140=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_140=1.27e-10
.param mcm2l1_cf_w_1_120_s_0_140=2.57e-12
.param mcm2l1_ca_w_1_120_s_0_175=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_175=1.22e-10
.param mcm2l1_cf_w_1_120_s_0_175=3.21e-12
.param mcm2l1_ca_w_1_120_s_0_210=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_210=1.16e-10
.param mcm2l1_cf_w_1_120_s_0_210=3.85e-12
.param mcm2l1_ca_w_1_120_s_0_280=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_280=1.02e-10
.param mcm2l1_cf_w_1_120_s_0_280=5.10e-12
.param mcm2l1_ca_w_1_120_s_0_350=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_350=8.96e-11
.param mcm2l1_cf_w_1_120_s_0_350=6.32e-12
.param mcm2l1_ca_w_1_120_s_0_420=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_420=7.92e-11
.param mcm2l1_cf_w_1_120_s_0_420=7.52e-12
.param mcm2l1_ca_w_1_120_s_0_560=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_560=6.41e-11
.param mcm2l1_cf_w_1_120_s_0_560=9.79e-12
.param mcm2l1_ca_w_1_120_s_0_840=3.70e-05
.param mcm2l1_cc_w_1_120_s_0_840=4.73e-11
.param mcm2l1_cf_w_1_120_s_0_840=1.40e-11
.param mcm2l1_ca_w_1_120_s_1_540=3.70e-05
.param mcm2l1_cc_w_1_120_s_1_540=2.86e-11
.param mcm2l1_cf_w_1_120_s_1_540=2.25e-11
.param mcm2l1_ca_w_1_120_s_3_500=3.70e-05
.param mcm2l1_cc_w_1_120_s_3_500=1.18e-11
.param mcm2l1_cf_w_1_120_s_3_500=3.52e-11
.param mcm2m1_ca_w_0_140_s_0_140=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_140=9.46e-11
.param mcm2m1_cf_w_0_140_s_0_140=8.24e-12
.param mcm2m1_ca_w_0_140_s_0_175=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_175=9.27e-11
.param mcm2m1_cf_w_0_140_s_0_175=1.04e-11
.param mcm2m1_ca_w_0_140_s_0_210=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_210=8.69e-11
.param mcm2m1_cf_w_0_140_s_0_210=1.25e-11
.param mcm2m1_ca_w_0_140_s_0_280=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_280=7.48e-11
.param mcm2m1_cf_w_0_140_s_0_280=1.65e-11
.param mcm2m1_ca_w_0_140_s_0_350=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_350=6.32e-11
.param mcm2m1_cf_w_0_140_s_0_350=2.01e-11
.param mcm2m1_ca_w_0_140_s_0_420=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_420=5.31e-11
.param mcm2m1_cf_w_0_140_s_0_420=2.34e-11
.param mcm2m1_ca_w_0_140_s_0_560=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_560=4.01e-11
.param mcm2m1_cf_w_0_140_s_0_560=2.91e-11
.param mcm2m1_ca_w_0_140_s_0_840=1.28e-04
.param mcm2m1_cc_w_0_140_s_0_840=2.60e-11
.param mcm2m1_cf_w_0_140_s_0_840=3.77e-11
.param mcm2m1_ca_w_0_140_s_1_540=1.28e-04
.param mcm2m1_cc_w_0_140_s_1_540=1.19e-11
.param mcm2m1_cf_w_0_140_s_1_540=4.94e-11
.param mcm2m1_ca_w_0_140_s_3_500=1.28e-04
.param mcm2m1_cc_w_0_140_s_3_500=3.35e-12
.param mcm2m1_cf_w_0_140_s_3_500=5.79e-11
.param mcm2m1_ca_w_1_120_s_0_140=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_140=1.13e-10
.param mcm2m1_cf_w_1_120_s_0_140=8.25e-12
.param mcm2m1_ca_w_1_120_s_0_175=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_175=1.09e-10
.param mcm2m1_cf_w_1_120_s_0_175=1.05e-11
.param mcm2m1_ca_w_1_120_s_0_210=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_210=1.02e-10
.param mcm2m1_cf_w_1_120_s_0_210=1.25e-11
.param mcm2m1_ca_w_1_120_s_0_280=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_280=8.91e-11
.param mcm2m1_cf_w_1_120_s_0_280=1.65e-11
.param mcm2m1_ca_w_1_120_s_0_350=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_350=7.62e-11
.param mcm2m1_cf_w_1_120_s_0_350=2.01e-11
.param mcm2m1_ca_w_1_120_s_0_420=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_420=6.60e-11
.param mcm2m1_cf_w_1_120_s_0_420=2.34e-11
.param mcm2m1_ca_w_1_120_s_0_560=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_560=5.15e-11
.param mcm2m1_cf_w_1_120_s_0_560=2.91e-11
.param mcm2m1_ca_w_1_120_s_0_840=1.28e-04
.param mcm2m1_cc_w_1_120_s_0_840=3.55e-11
.param mcm2m1_cf_w_1_120_s_0_840=3.78e-11
.param mcm2m1_ca_w_1_120_s_1_540=1.28e-04
.param mcm2m1_cc_w_1_120_s_1_540=1.90e-11
.param mcm2m1_cf_w_1_120_s_1_540=5.05e-11
.param mcm2m1_ca_w_1_120_s_3_500=1.28e-04
.param mcm2m1_cc_w_1_120_s_3_500=6.75e-12
.param mcm2m1_cf_w_1_120_s_3_500=6.23e-11
.param mcm3f_ca_w_0_300_s_0_300=1.26e-05
.param mcm3f_cc_w_0_300_s_0_300=1.06e-10
.param mcm3f_cf_w_0_300_s_0_300=1.86e-12
.param mcm3f_ca_w_0_300_s_0_360=1.26e-05
.param mcm3f_cc_w_0_300_s_0_360=9.95e-11
.param mcm3f_cf_w_0_300_s_0_360=2.22e-12
.param mcm3f_ca_w_0_300_s_0_450=1.26e-05
.param mcm3f_cc_w_0_300_s_0_450=8.98e-11
.param mcm3f_cf_w_0_300_s_0_450=2.79e-12
.param mcm3f_ca_w_0_300_s_0_600=1.26e-05
.param mcm3f_cc_w_0_300_s_0_600=7.73e-11
.param mcm3f_cf_w_0_300_s_0_600=3.70e-12
.param mcm3f_ca_w_0_300_s_0_800=1.26e-05
.param mcm3f_cc_w_0_300_s_0_800=6.53e-11
.param mcm3f_cf_w_0_300_s_0_800=4.80e-12
.param mcm3f_ca_w_0_300_s_1_000=1.26e-05
.param mcm3f_cc_w_0_300_s_1_000=5.62e-11
.param mcm3f_cf_w_0_300_s_1_000=5.93e-12
.param mcm3f_ca_w_0_300_s_1_200=1.26e-05
.param mcm3f_cc_w_0_300_s_1_200=4.95e-11
.param mcm3f_cf_w_0_300_s_1_200=7.00e-12
.param mcm3f_ca_w_0_300_s_2_100=1.26e-05
.param mcm3f_cc_w_0_300_s_2_100=3.26e-11
.param mcm3f_cf_w_0_300_s_2_100=1.18e-11
.param mcm3f_ca_w_0_300_s_3_300=1.26e-05
.param mcm3f_cc_w_0_300_s_3_300=2.26e-11
.param mcm3f_cf_w_0_300_s_3_300=1.64e-11
.param mcm3f_ca_w_0_300_s_9_000=1.26e-05
.param mcm3f_cc_w_0_300_s_9_000=6.81e-12
.param mcm3f_cf_w_0_300_s_9_000=2.82e-11
.param mcm3f_ca_w_2_400_s_0_300=1.26e-05
.param mcm3f_cc_w_2_400_s_0_300=1.32e-10
.param mcm3f_cf_w_2_400_s_0_300=1.89e-12
.param mcm3f_ca_w_2_400_s_0_360=1.26e-05
.param mcm3f_cc_w_2_400_s_0_360=1.23e-10
.param mcm3f_cf_w_2_400_s_0_360=2.26e-12
.param mcm3f_ca_w_2_400_s_0_450=1.26e-05
.param mcm3f_cc_w_2_400_s_0_450=1.12e-10
.param mcm3f_cf_w_2_400_s_0_450=2.80e-12
.param mcm3f_ca_w_2_400_s_0_600=1.26e-05
.param mcm3f_cc_w_2_400_s_0_600=9.72e-11
.param mcm3f_cf_w_2_400_s_0_600=3.69e-12
.param mcm3f_ca_w_2_400_s_0_800=1.26e-05
.param mcm3f_cc_w_2_400_s_0_800=8.27e-11
.param mcm3f_cf_w_2_400_s_0_800=4.86e-12
.param mcm3f_ca_w_2_400_s_1_000=1.26e-05
.param mcm3f_cc_w_2_400_s_1_000=7.19e-11
.param mcm3f_cf_w_2_400_s_1_000=6.00e-12
.param mcm3f_ca_w_2_400_s_1_200=1.26e-05
.param mcm3f_cc_w_2_400_s_1_200=6.38e-11
.param mcm3f_cf_w_2_400_s_1_200=7.11e-12
.param mcm3f_ca_w_2_400_s_2_100=1.26e-05
.param mcm3f_cc_w_2_400_s_2_100=4.35e-11
.param mcm3f_cf_w_2_400_s_2_100=1.17e-11
.param mcm3f_ca_w_2_400_s_3_300=1.26e-05
.param mcm3f_cc_w_2_400_s_3_300=3.06e-11
.param mcm3f_cf_w_2_400_s_3_300=1.69e-11
.param mcm3f_ca_w_2_400_s_9_000=1.26e-05
.param mcm3f_cc_w_2_400_s_9_000=1.05e-11
.param mcm3f_cf_w_2_400_s_9_000=3.09e-11
.param mcm3d_ca_w_0_300_s_0_300=1.42e-05
.param mcm3d_cc_w_0_300_s_0_300=1.06e-10
.param mcm3d_cf_w_0_300_s_0_300=2.09e-12
.param mcm3d_ca_w_0_300_s_0_360=1.42e-05
.param mcm3d_cc_w_0_300_s_0_360=9.90e-11
.param mcm3d_cf_w_0_300_s_0_360=2.50e-12
.param mcm3d_ca_w_0_300_s_0_450=1.42e-05
.param mcm3d_cc_w_0_300_s_0_450=8.93e-11
.param mcm3d_cf_w_0_300_s_0_450=3.13e-12
.param mcm3d_ca_w_0_300_s_0_600=1.42e-05
.param mcm3d_cc_w_0_300_s_0_600=7.68e-11
.param mcm3d_cf_w_0_300_s_0_600=4.15e-12
.param mcm3d_ca_w_0_300_s_0_800=1.42e-05
.param mcm3d_cc_w_0_300_s_0_800=6.46e-11
.param mcm3d_cf_w_0_300_s_0_800=5.39e-12
.param mcm3d_ca_w_0_300_s_1_000=1.42e-05
.param mcm3d_cc_w_0_300_s_1_000=5.55e-11
.param mcm3d_cf_w_0_300_s_1_000=6.64e-12
.param mcm3d_ca_w_0_300_s_1_200=1.42e-05
.param mcm3d_cc_w_0_300_s_1_200=4.86e-11
.param mcm3d_cf_w_0_300_s_1_200=7.84e-12
.param mcm3d_ca_w_0_300_s_2_100=1.42e-05
.param mcm3d_cc_w_0_300_s_2_100=3.16e-11
.param mcm3d_cf_w_0_300_s_2_100=1.31e-11
.param mcm3d_ca_w_0_300_s_3_300=1.42e-05
.param mcm3d_cc_w_0_300_s_3_300=2.16e-11
.param mcm3d_cf_w_0_300_s_3_300=1.80e-11
.param mcm3d_ca_w_0_300_s_9_000=1.42e-05
.param mcm3d_cc_w_0_300_s_9_000=6.17e-12
.param mcm3d_cf_w_0_300_s_9_000=2.99e-11
.param mcm3d_ca_w_2_400_s_0_300=1.42e-05
.param mcm3d_cc_w_2_400_s_0_300=1.30e-10
.param mcm3d_cf_w_2_400_s_0_300=2.14e-12
.param mcm3d_ca_w_2_400_s_0_360=1.42e-05
.param mcm3d_cc_w_2_400_s_0_360=1.22e-10
.param mcm3d_cf_w_2_400_s_0_360=2.55e-12
.param mcm3d_ca_w_2_400_s_0_450=1.42e-05
.param mcm3d_cc_w_2_400_s_0_450=1.11e-10
.param mcm3d_cf_w_2_400_s_0_450=3.16e-12
.param mcm3d_ca_w_2_400_s_0_600=1.42e-05
.param mcm3d_cc_w_2_400_s_0_600=9.60e-11
.param mcm3d_cf_w_2_400_s_0_600=4.15e-12
.param mcm3d_ca_w_2_400_s_0_800=1.42e-05
.param mcm3d_cc_w_2_400_s_0_800=8.14e-11
.param mcm3d_cf_w_2_400_s_0_800=5.45e-12
.param mcm3d_ca_w_2_400_s_1_000=1.42e-05
.param mcm3d_cc_w_2_400_s_1_000=7.06e-11
.param mcm3d_cf_w_2_400_s_1_000=6.72e-12
.param mcm3d_ca_w_2_400_s_1_200=1.42e-05
.param mcm3d_cc_w_2_400_s_1_200=6.25e-11
.param mcm3d_cf_w_2_400_s_1_200=7.94e-12
.param mcm3d_ca_w_2_400_s_2_100=1.42e-05
.param mcm3d_cc_w_2_400_s_2_100=4.22e-11
.param mcm3d_cf_w_2_400_s_2_100=1.30e-11
.param mcm3d_ca_w_2_400_s_3_300=1.42e-05
.param mcm3d_cc_w_2_400_s_3_300=2.95e-11
.param mcm3d_cf_w_2_400_s_3_300=1.86e-11
.param mcm3d_ca_w_2_400_s_9_000=1.42e-05
.param mcm3d_cc_w_2_400_s_9_000=9.73e-12
.param mcm3d_cf_w_2_400_s_9_000=3.28e-11
.param mcm3p1_ca_w_0_300_s_0_300=1.58e-05
.param mcm3p1_cc_w_0_300_s_0_300=1.06e-10
.param mcm3p1_cf_w_0_300_s_0_300=2.34e-12
.param mcm3p1_ca_w_0_300_s_0_360=1.58e-05
.param mcm3p1_cc_w_0_300_s_0_360=9.84e-11
.param mcm3p1_cf_w_0_300_s_0_360=2.80e-12
.param mcm3p1_ca_w_0_300_s_0_450=1.58e-05
.param mcm3p1_cc_w_0_300_s_0_450=8.89e-11
.param mcm3p1_cf_w_0_300_s_0_450=3.50e-12
.param mcm3p1_ca_w_0_300_s_0_600=1.58e-05
.param mcm3p1_cc_w_0_300_s_0_600=7.62e-11
.param mcm3p1_cf_w_0_300_s_0_600=4.63e-12
.param mcm3p1_ca_w_0_300_s_0_800=1.58e-05
.param mcm3p1_cc_w_0_300_s_0_800=6.40e-11
.param mcm3p1_cf_w_0_300_s_0_800=6.00e-12
.param mcm3p1_ca_w_0_300_s_1_000=1.58e-05
.param mcm3p1_cc_w_0_300_s_1_000=5.48e-11
.param mcm3p1_cf_w_0_300_s_1_000=7.39e-12
.param mcm3p1_ca_w_0_300_s_1_200=1.58e-05
.param mcm3p1_cc_w_0_300_s_1_200=4.79e-11
.param mcm3p1_cf_w_0_300_s_1_200=8.70e-12
.param mcm3p1_ca_w_0_300_s_2_100=1.58e-05
.param mcm3p1_cc_w_0_300_s_2_100=3.07e-11
.param mcm3p1_cf_w_0_300_s_2_100=1.44e-11
.param mcm3p1_ca_w_0_300_s_3_300=1.58e-05
.param mcm3p1_cc_w_0_300_s_3_300=2.06e-11
.param mcm3p1_cf_w_0_300_s_3_300=1.96e-11
.param mcm3p1_ca_w_0_300_s_9_000=1.58e-05
.param mcm3p1_cc_w_0_300_s_9_000=5.69e-12
.param mcm3p1_cf_w_0_300_s_9_000=3.15e-11
.param mcm3p1_ca_w_2_400_s_0_300=1.58e-05
.param mcm3p1_cc_w_2_400_s_0_300=1.29e-10
.param mcm3p1_cf_w_2_400_s_0_300=2.42e-12
.param mcm3p1_ca_w_2_400_s_0_360=1.58e-05
.param mcm3p1_cc_w_2_400_s_0_360=1.21e-10
.param mcm3p1_cf_w_2_400_s_0_360=2.87e-12
.param mcm3p1_ca_w_2_400_s_0_450=1.58e-05
.param mcm3p1_cc_w_2_400_s_0_450=1.09e-10
.param mcm3p1_cf_w_2_400_s_0_450=3.55e-12
.param mcm3p1_ca_w_2_400_s_0_600=1.58e-05
.param mcm3p1_cc_w_2_400_s_0_600=9.49e-11
.param mcm3p1_cf_w_2_400_s_0_600=4.66e-12
.param mcm3p1_ca_w_2_400_s_0_800=1.58e-05
.param mcm3p1_cc_w_2_400_s_0_800=8.02e-11
.param mcm3p1_cf_w_2_400_s_0_800=6.10e-12
.param mcm3p1_ca_w_2_400_s_1_000=1.58e-05
.param mcm3p1_cc_w_2_400_s_1_000=6.94e-11
.param mcm3p1_cf_w_2_400_s_1_000=7.49e-12
.param mcm3p1_ca_w_2_400_s_1_200=1.58e-05
.param mcm3p1_cc_w_2_400_s_1_200=6.13e-11
.param mcm3p1_cf_w_2_400_s_1_200=8.85e-12
.param mcm3p1_ca_w_2_400_s_2_100=1.58e-05
.param mcm3p1_cc_w_2_400_s_2_100=4.10e-11
.param mcm3p1_cf_w_2_400_s_2_100=1.43e-11
.param mcm3p1_ca_w_2_400_s_3_300=1.58e-05
.param mcm3p1_cc_w_2_400_s_3_300=2.83e-11
.param mcm3p1_cf_w_2_400_s_3_300=2.03e-11
.param mcm3p1_ca_w_2_400_s_9_000=1.58e-05
.param mcm3p1_cc_w_2_400_s_9_000=9.05e-12
.param mcm3p1_cf_w_2_400_s_9_000=3.46e-11
.param mcm3l1_ca_w_0_300_s_0_300=2.02e-05
.param mcm3l1_cc_w_0_300_s_0_300=1.05e-10
.param mcm3l1_cf_w_0_300_s_0_300=2.95e-12
.param mcm3l1_ca_w_0_300_s_0_360=2.02e-05
.param mcm3l1_cc_w_0_300_s_0_360=9.73e-11
.param mcm3l1_cf_w_0_300_s_0_360=3.52e-12
.param mcm3l1_ca_w_0_300_s_0_450=2.02e-05
.param mcm3l1_cc_w_0_300_s_0_450=8.75e-11
.param mcm3l1_cf_w_0_300_s_0_450=4.38e-12
.param mcm3l1_ca_w_0_300_s_0_600=2.02e-05
.param mcm3l1_cc_w_0_300_s_0_600=7.49e-11
.param mcm3l1_cf_w_0_300_s_0_600=5.78e-12
.param mcm3l1_ca_w_0_300_s_0_800=2.02e-05
.param mcm3l1_cc_w_0_300_s_0_800=6.24e-11
.param mcm3l1_cf_w_0_300_s_0_800=7.48e-12
.param mcm3l1_ca_w_0_300_s_1_000=2.02e-05
.param mcm3l1_cc_w_0_300_s_1_000=5.32e-11
.param mcm3l1_cf_w_0_300_s_1_000=9.16e-12
.param mcm3l1_ca_w_0_300_s_1_200=2.02e-05
.param mcm3l1_cc_w_0_300_s_1_200=4.62e-11
.param mcm3l1_cf_w_0_300_s_1_200=1.08e-11
.param mcm3l1_ca_w_0_300_s_2_100=2.02e-05
.param mcm3l1_cc_w_0_300_s_2_100=2.86e-11
.param mcm3l1_cf_w_0_300_s_2_100=1.74e-11
.param mcm3l1_ca_w_0_300_s_3_300=2.02e-05
.param mcm3l1_cc_w_0_300_s_3_300=1.86e-11
.param mcm3l1_cf_w_0_300_s_3_300=2.32e-11
.param mcm3l1_ca_w_0_300_s_9_000=2.02e-05
.param mcm3l1_cc_w_0_300_s_9_000=4.69e-12
.param mcm3l1_cf_w_0_300_s_9_000=3.48e-11
.param mcm3l1_ca_w_2_400_s_0_300=2.02e-05
.param mcm3l1_cc_w_2_400_s_0_300=1.27e-10
.param mcm3l1_cf_w_2_400_s_0_300=2.99e-12
.param mcm3l1_ca_w_2_400_s_0_360=2.02e-05
.param mcm3l1_cc_w_2_400_s_0_360=1.18e-10
.param mcm3l1_cf_w_2_400_s_0_360=3.56e-12
.param mcm3l1_ca_w_2_400_s_0_450=2.02e-05
.param mcm3l1_cc_w_2_400_s_0_450=1.07e-10
.param mcm3l1_cf_w_2_400_s_0_450=4.41e-12
.param mcm3l1_ca_w_2_400_s_0_600=2.02e-05
.param mcm3l1_cc_w_2_400_s_0_600=9.24e-11
.param mcm3l1_cf_w_2_400_s_0_600=5.78e-12
.param mcm3l1_ca_w_2_400_s_0_800=2.02e-05
.param mcm3l1_cc_w_2_400_s_0_800=7.77e-11
.param mcm3l1_cf_w_2_400_s_0_800=7.55e-12
.param mcm3l1_ca_w_2_400_s_1_000=2.02e-05
.param mcm3l1_cc_w_2_400_s_1_000=6.68e-11
.param mcm3l1_cf_w_2_400_s_1_000=9.25e-12
.param mcm3l1_ca_w_2_400_s_1_200=2.02e-05
.param mcm3l1_cc_w_2_400_s_1_200=5.87e-11
.param mcm3l1_cf_w_2_400_s_1_200=1.09e-11
.param mcm3l1_ca_w_2_400_s_2_100=2.02e-05
.param mcm3l1_cc_w_2_400_s_2_100=3.86e-11
.param mcm3l1_cf_w_2_400_s_2_100=1.73e-11
.param mcm3l1_ca_w_2_400_s_3_300=2.02e-05
.param mcm3l1_cc_w_2_400_s_3_300=2.60e-11
.param mcm3l1_cf_w_2_400_s_3_300=2.40e-11
.param mcm3l1_ca_w_2_400_s_9_000=2.02e-05
.param mcm3l1_cc_w_2_400_s_9_000=7.85e-12
.param mcm3l1_cf_w_2_400_s_9_000=3.84e-11
.param mcm3m1_ca_w_0_300_s_0_300=3.29e-05
.param mcm3m1_cc_w_0_300_s_0_300=1.02e-10
.param mcm3m1_cf_w_0_300_s_0_300=4.72e-12
.param mcm3m1_ca_w_0_300_s_0_360=3.29e-05
.param mcm3m1_cc_w_0_300_s_0_360=9.42e-11
.param mcm3m1_cf_w_0_300_s_0_360=5.62e-12
.param mcm3m1_ca_w_0_300_s_0_450=3.29e-05
.param mcm3m1_cc_w_0_300_s_0_450=8.43e-11
.param mcm3m1_cf_w_0_300_s_0_450=6.94e-12
.param mcm3m1_ca_w_0_300_s_0_600=3.29e-05
.param mcm3m1_cc_w_0_300_s_0_600=7.13e-11
.param mcm3m1_cf_w_0_300_s_0_600=9.07e-12
.param mcm3m1_ca_w_0_300_s_0_800=3.29e-05
.param mcm3m1_cc_w_0_300_s_0_800=5.87e-11
.param mcm3m1_cf_w_0_300_s_0_800=1.16e-11
.param mcm3m1_ca_w_0_300_s_1_000=3.29e-05
.param mcm3m1_cc_w_0_300_s_1_000=4.91e-11
.param mcm3m1_cf_w_0_300_s_1_000=1.41e-11
.param mcm3m1_ca_w_0_300_s_1_200=3.29e-05
.param mcm3m1_cc_w_0_300_s_1_200=4.20e-11
.param mcm3m1_cf_w_0_300_s_1_200=1.64e-11
.param mcm3m1_ca_w_0_300_s_2_100=3.29e-05
.param mcm3m1_cc_w_0_300_s_2_100=2.43e-11
.param mcm3m1_cf_w_0_300_s_2_100=2.51e-11
.param mcm3m1_ca_w_0_300_s_3_300=3.29e-05
.param mcm3m1_cc_w_0_300_s_3_300=1.48e-11
.param mcm3m1_cf_w_0_300_s_3_300=3.17e-11
.param mcm3m1_ca_w_0_300_s_9_000=3.29e-05
.param mcm3m1_cc_w_0_300_s_9_000=3.27e-12
.param mcm3m1_cf_w_0_300_s_9_000=4.21e-11
.param mcm3m1_ca_w_2_400_s_0_300=3.29e-05
.param mcm3m1_cc_w_2_400_s_0_300=1.21e-10
.param mcm3m1_cf_w_2_400_s_0_300=4.73e-12
.param mcm3m1_ca_w_2_400_s_0_360=3.29e-05
.param mcm3m1_cc_w_2_400_s_0_360=1.13e-10
.param mcm3m1_cf_w_2_400_s_0_360=5.64e-12
.param mcm3m1_ca_w_2_400_s_0_450=3.29e-05
.param mcm3m1_cc_w_2_400_s_0_450=1.02e-10
.param mcm3m1_cf_w_2_400_s_0_450=6.95e-12
.param mcm3m1_ca_w_2_400_s_0_600=3.29e-05
.param mcm3m1_cc_w_2_400_s_0_600=8.70e-11
.param mcm3m1_cf_w_2_400_s_0_600=9.05e-12
.param mcm3m1_ca_w_2_400_s_0_800=3.29e-05
.param mcm3m1_cc_w_2_400_s_0_800=7.25e-11
.param mcm3m1_cf_w_2_400_s_0_800=1.17e-11
.param mcm3m1_ca_w_2_400_s_1_000=3.29e-05
.param mcm3m1_cc_w_2_400_s_1_000=6.18e-11
.param mcm3m1_cf_w_2_400_s_1_000=1.42e-11
.param mcm3m1_ca_w_2_400_s_1_200=3.29e-05
.param mcm3m1_cc_w_2_400_s_1_200=5.38e-11
.param mcm3m1_cf_w_2_400_s_1_200=1.65e-11
.param mcm3m1_ca_w_2_400_s_2_100=3.29e-05
.param mcm3m1_cc_w_2_400_s_2_100=3.39e-11
.param mcm3m1_cf_w_2_400_s_2_100=2.49e-11
.param mcm3m1_ca_w_2_400_s_3_300=3.29e-05
.param mcm3m1_cc_w_2_400_s_3_300=2.20e-11
.param mcm3m1_cf_w_2_400_s_3_300=3.27e-11
.param mcm3m1_ca_w_2_400_s_9_000=3.29e-05
.param mcm3m1_cc_w_2_400_s_9_000=6.00e-12
.param mcm3m1_cf_w_2_400_s_9_000=4.65e-11
.param mcm3m2_ca_w_0_300_s_0_300=8.22e-05
.param mcm3m2_cc_w_0_300_s_0_300=9.39e-11
.param mcm3m2_cf_w_0_300_s_0_300=1.11e-11
.param mcm3m2_ca_w_0_300_s_0_360=8.22e-05
.param mcm3m2_cc_w_0_300_s_0_360=8.63e-11
.param mcm3m2_cf_w_0_300_s_0_360=1.30e-11
.param mcm3m2_ca_w_0_300_s_0_450=8.22e-05
.param mcm3m2_cc_w_0_300_s_0_450=7.63e-11
.param mcm3m2_cf_w_0_300_s_0_450=1.57e-11
.param mcm3m2_ca_w_0_300_s_0_600=8.22e-05
.param mcm3m2_cc_w_0_300_s_0_600=6.30e-11
.param mcm3m2_cf_w_0_300_s_0_600=1.99e-11
.param mcm3m2_ca_w_0_300_s_0_800=8.22e-05
.param mcm3m2_cc_w_0_300_s_0_800=5.03e-11
.param mcm3m2_cf_w_0_300_s_0_800=2.45e-11
.param mcm3m2_ca_w_0_300_s_1_000=8.22e-05
.param mcm3m2_cc_w_0_300_s_1_000=4.10e-11
.param mcm3m2_cf_w_0_300_s_1_000=2.85e-11
.param mcm3m2_ca_w_0_300_s_1_200=8.22e-05
.param mcm3m2_cc_w_0_300_s_1_200=3.42e-11
.param mcm3m2_cf_w_0_300_s_1_200=3.19e-11
.param mcm3m2_ca_w_0_300_s_2_100=8.22e-05
.param mcm3m2_cc_w_0_300_s_2_100=1.76e-11
.param mcm3m2_cf_w_0_300_s_2_100=4.31e-11
.param mcm3m2_ca_w_0_300_s_3_300=8.22e-05
.param mcm3m2_cc_w_0_300_s_3_300=9.90e-12
.param mcm3m2_cf_w_0_300_s_3_300=4.95e-11
.param mcm3m2_ca_w_0_300_s_9_000=8.22e-05
.param mcm3m2_cc_w_0_300_s_9_000=1.95e-12
.param mcm3m2_cf_w_0_300_s_9_000=5.72e-11
.param mcm3m2_ca_w_2_400_s_0_300=8.22e-05
.param mcm3m2_cc_w_2_400_s_0_300=1.11e-10
.param mcm3m2_cf_w_2_400_s_0_300=1.11e-11
.param mcm3m2_ca_w_2_400_s_0_360=8.22e-05
.param mcm3m2_cc_w_2_400_s_0_360=1.03e-10
.param mcm3m2_cf_w_2_400_s_0_360=1.30e-11
.param mcm3m2_ca_w_2_400_s_0_450=8.22e-05
.param mcm3m2_cc_w_2_400_s_0_450=9.20e-11
.param mcm3m2_cf_w_2_400_s_0_450=1.57e-11
.param mcm3m2_ca_w_2_400_s_0_600=8.22e-05
.param mcm3m2_cc_w_2_400_s_0_600=7.76e-11
.param mcm3m2_cf_w_2_400_s_0_600=1.98e-11
.param mcm3m2_ca_w_2_400_s_0_800=8.22e-05
.param mcm3m2_cc_w_2_400_s_0_800=6.33e-11
.param mcm3m2_cf_w_2_400_s_0_800=2.45e-11
.param mcm3m2_ca_w_2_400_s_1_000=8.22e-05
.param mcm3m2_cc_w_2_400_s_1_000=5.31e-11
.param mcm3m2_cf_w_2_400_s_1_000=2.86e-11
.param mcm3m2_ca_w_2_400_s_1_200=8.22e-05
.param mcm3m2_cc_w_2_400_s_1_200=4.56e-11
.param mcm3m2_cf_w_2_400_s_1_200=3.20e-11
.param mcm3m2_ca_w_2_400_s_2_100=8.22e-05
.param mcm3m2_cc_w_2_400_s_2_100=2.72e-11
.param mcm3m2_cf_w_2_400_s_2_100=4.29e-11
.param mcm3m2_ca_w_2_400_s_3_300=8.22e-05
.param mcm3m2_cc_w_2_400_s_3_300=1.68e-11
.param mcm3m2_cf_w_2_400_s_3_300=5.12e-11
.param mcm3m2_ca_w_2_400_s_9_000=8.22e-05
.param mcm3m2_cc_w_2_400_s_9_000=4.25e-12
.param mcm3m2_cf_w_2_400_s_9_000=6.29e-11
.param mcm4f_ca_w_0_300_s_0_300=8.67e-06
.param mcm4f_cc_w_0_300_s_0_300=1.08e-10
.param mcm4f_cf_w_0_300_s_0_300=1.29e-12
.param mcm4f_ca_w_0_300_s_0_360=8.67e-06
.param mcm4f_cc_w_0_300_s_0_360=1.01e-10
.param mcm4f_cf_w_0_300_s_0_360=1.54e-12
.param mcm4f_ca_w_0_300_s_0_450=8.67e-06
.param mcm4f_cc_w_0_300_s_0_450=9.17e-11
.param mcm4f_cf_w_0_300_s_0_450=1.94e-12
.param mcm4f_ca_w_0_300_s_0_600=8.67e-06
.param mcm4f_cc_w_0_300_s_0_600=7.96e-11
.param mcm4f_cf_w_0_300_s_0_600=2.59e-12
.param mcm4f_ca_w_0_300_s_0_800=8.67e-06
.param mcm4f_cc_w_0_300_s_0_800=6.78e-11
.param mcm4f_cf_w_0_300_s_0_800=3.35e-12
.param mcm4f_ca_w_0_300_s_1_000=8.67e-06
.param mcm4f_cc_w_0_300_s_1_000=5.90e-11
.param mcm4f_cf_w_0_300_s_1_000=4.16e-12
.param mcm4f_ca_w_0_300_s_1_200=8.67e-06
.param mcm4f_cc_w_0_300_s_1_200=5.24e-11
.param mcm4f_cf_w_0_300_s_1_200=4.94e-12
.param mcm4f_ca_w_0_300_s_2_100=8.67e-06
.param mcm4f_cc_w_0_300_s_2_100=3.60e-11
.param mcm4f_cf_w_0_300_s_2_100=8.49e-12
.param mcm4f_ca_w_0_300_s_3_300=8.67e-06
.param mcm4f_cc_w_0_300_s_3_300=2.59e-11
.param mcm4f_cf_w_0_300_s_3_300=1.21e-11
.param mcm4f_ca_w_0_300_s_9_000=8.67e-06
.param mcm4f_cc_w_0_300_s_9_000=8.98e-12
.param mcm4f_cf_w_0_300_s_9_000=2.31e-11
.param mcm4f_ca_w_2_400_s_0_300=8.67e-06
.param mcm4f_cc_w_2_400_s_0_300=1.36e-10
.param mcm4f_cf_w_2_400_s_0_300=1.31e-12
.param mcm4f_ca_w_2_400_s_0_360=8.67e-06
.param mcm4f_cc_w_2_400_s_0_360=1.28e-10
.param mcm4f_cf_w_2_400_s_0_360=1.56e-12
.param mcm4f_ca_w_2_400_s_0_450=8.67e-06
.param mcm4f_cc_w_2_400_s_0_450=1.17e-10
.param mcm4f_cf_w_2_400_s_0_450=1.94e-12
.param mcm4f_ca_w_2_400_s_0_600=8.67e-06
.param mcm4f_cc_w_2_400_s_0_600=1.02e-10
.param mcm4f_cf_w_2_400_s_0_600=2.57e-12
.param mcm4f_ca_w_2_400_s_0_800=8.67e-06
.param mcm4f_cc_w_2_400_s_0_800=8.75e-11
.param mcm4f_cf_w_2_400_s_0_800=3.39e-12
.param mcm4f_ca_w_2_400_s_1_000=8.67e-06
.param mcm4f_cc_w_2_400_s_1_000=7.66e-11
.param mcm4f_cf_w_2_400_s_1_000=4.20e-12
.param mcm4f_ca_w_2_400_s_1_200=8.67e-06
.param mcm4f_cc_w_2_400_s_1_200=6.84e-11
.param mcm4f_cf_w_2_400_s_1_200=4.99e-12
.param mcm4f_ca_w_2_400_s_2_100=8.67e-06
.param mcm4f_cc_w_2_400_s_2_100=4.77e-11
.param mcm4f_cf_w_2_400_s_2_100=8.38e-12
.param mcm4f_ca_w_2_400_s_3_300=8.67e-06
.param mcm4f_cc_w_2_400_s_3_300=3.44e-11
.param mcm4f_cf_w_2_400_s_3_300=1.24e-11
.param mcm4f_ca_w_2_400_s_9_000=8.67e-06
.param mcm4f_cc_w_2_400_s_9_000=1.29e-11
.param mcm4f_cf_w_2_400_s_9_000=2.51e-11
.param mcm4d_ca_w_0_300_s_0_300=9.41e-06
.param mcm4d_cc_w_0_300_s_0_300=1.08e-10
.param mcm4d_cf_w_0_300_s_0_300=1.39e-12
.param mcm4d_ca_w_0_300_s_0_360=9.41e-06
.param mcm4d_cc_w_0_300_s_0_360=1.01e-10
.param mcm4d_cf_w_0_300_s_0_360=1.67e-12
.param mcm4d_ca_w_0_300_s_0_450=9.41e-06
.param mcm4d_cc_w_0_300_s_0_450=9.14e-11
.param mcm4d_cf_w_0_300_s_0_450=2.10e-12
.param mcm4d_ca_w_0_300_s_0_600=9.41e-06
.param mcm4d_cc_w_0_300_s_0_600=7.93e-11
.param mcm4d_cf_w_0_300_s_0_600=2.80e-12
.param mcm4d_ca_w_0_300_s_0_800=9.41e-06
.param mcm4d_cc_w_0_300_s_0_800=6.75e-11
.param mcm4d_cf_w_0_300_s_0_800=3.63e-12
.param mcm4d_ca_w_0_300_s_1_000=9.41e-06
.param mcm4d_cc_w_0_300_s_1_000=5.87e-11
.param mcm4d_cf_w_0_300_s_1_000=4.49e-12
.param mcm4d_ca_w_0_300_s_1_200=9.41e-06
.param mcm4d_cc_w_0_300_s_1_200=5.20e-11
.param mcm4d_cf_w_0_300_s_1_200=5.34e-12
.param mcm4d_ca_w_0_300_s_2_100=9.41e-06
.param mcm4d_cc_w_0_300_s_2_100=3.54e-11
.param mcm4d_cf_w_0_300_s_2_100=9.13e-12
.param mcm4d_ca_w_0_300_s_3_300=9.41e-06
.param mcm4d_cc_w_0_300_s_3_300=2.53e-11
.param mcm4d_cf_w_0_300_s_3_300=1.29e-11
.param mcm4d_ca_w_0_300_s_9_000=9.41e-06
.param mcm4d_cc_w_0_300_s_9_000=8.44e-12
.param mcm4d_cf_w_0_300_s_9_000=2.42e-11
.param mcm4d_ca_w_2_400_s_0_300=9.41e-06
.param mcm4d_cc_w_2_400_s_0_300=1.36e-10
.param mcm4d_cf_w_2_400_s_0_300=1.42e-12
.param mcm4d_ca_w_2_400_s_0_360=9.41e-06
.param mcm4d_cc_w_2_400_s_0_360=1.27e-10
.param mcm4d_cf_w_2_400_s_0_360=1.69e-12
.param mcm4d_ca_w_2_400_s_0_450=9.41e-06
.param mcm4d_cc_w_2_400_s_0_450=1.17e-10
.param mcm4d_cf_w_2_400_s_0_450=2.10e-12
.param mcm4d_ca_w_2_400_s_0_600=9.41e-06
.param mcm4d_cc_w_2_400_s_0_600=1.01e-10
.param mcm4d_cf_w_2_400_s_0_600=2.78e-12
.param mcm4d_ca_w_2_400_s_0_800=9.41e-06
.param mcm4d_cc_w_2_400_s_0_800=8.67e-11
.param mcm4d_cf_w_2_400_s_0_800=3.67e-12
.param mcm4d_ca_w_2_400_s_1_000=9.41e-06
.param mcm4d_cc_w_2_400_s_1_000=7.59e-11
.param mcm4d_cf_w_2_400_s_1_000=4.54e-12
.param mcm4d_ca_w_2_400_s_1_200=9.41e-06
.param mcm4d_cc_w_2_400_s_1_200=6.77e-11
.param mcm4d_cf_w_2_400_s_1_200=5.40e-12
.param mcm4d_ca_w_2_400_s_2_100=9.41e-06
.param mcm4d_cc_w_2_400_s_2_100=4.69e-11
.param mcm4d_cf_w_2_400_s_2_100=9.02e-12
.param mcm4d_ca_w_2_400_s_3_300=9.41e-06
.param mcm4d_cc_w_2_400_s_3_300=3.36e-11
.param mcm4d_cf_w_2_400_s_3_300=1.33e-11
.param mcm4d_ca_w_2_400_s_9_000=9.41e-06
.param mcm4d_cc_w_2_400_s_9_000=1.23e-11
.param mcm4d_cf_w_2_400_s_9_000=2.63e-11
.param mcm4p1_ca_w_0_300_s_0_300=1.01e-05
.param mcm4p1_cc_w_0_300_s_0_300=1.07e-10
.param mcm4p1_cf_w_0_300_s_0_300=1.50e-12
.param mcm4p1_ca_w_0_300_s_0_360=1.01e-05
.param mcm4p1_cc_w_0_300_s_0_360=1.01e-10
.param mcm4p1_cf_w_0_300_s_0_360=1.80e-12
.param mcm4p1_ca_w_0_300_s_0_450=1.01e-05
.param mcm4p1_cc_w_0_300_s_0_450=9.12e-11
.param mcm4p1_cf_w_0_300_s_0_450=2.26e-12
.param mcm4p1_ca_w_0_300_s_0_600=1.01e-05
.param mcm4p1_cc_w_0_300_s_0_600=7.90e-11
.param mcm4p1_cf_w_0_300_s_0_600=3.01e-12
.param mcm4p1_ca_w_0_300_s_0_800=1.01e-05
.param mcm4p1_cc_w_0_300_s_0_800=6.71e-11
.param mcm4p1_cf_w_0_300_s_0_800=3.90e-12
.param mcm4p1_ca_w_0_300_s_1_000=1.01e-05
.param mcm4p1_cc_w_0_300_s_1_000=5.83e-11
.param mcm4p1_cf_w_0_300_s_1_000=4.83e-12
.param mcm4p1_ca_w_0_300_s_1_200=1.01e-05
.param mcm4p1_cc_w_0_300_s_1_200=5.16e-11
.param mcm4p1_cf_w_0_300_s_1_200=5.73e-12
.param mcm4p1_ca_w_0_300_s_2_100=1.01e-05
.param mcm4p1_cc_w_0_300_s_2_100=3.49e-11
.param mcm4p1_cf_w_0_300_s_2_100=9.75e-12
.param mcm4p1_ca_w_0_300_s_3_300=1.01e-05
.param mcm4p1_cc_w_0_300_s_3_300=2.47e-11
.param mcm4p1_cf_w_0_300_s_3_300=1.38e-11
.param mcm4p1_ca_w_0_300_s_9_000=1.01e-05
.param mcm4p1_cc_w_0_300_s_9_000=7.99e-12
.param mcm4p1_cf_w_0_300_s_9_000=2.53e-11
.param mcm4p1_ca_w_2_400_s_0_300=1.01e-05
.param mcm4p1_cc_w_2_400_s_0_300=1.35e-10
.param mcm4p1_cf_w_2_400_s_0_300=1.54e-12
.param mcm4p1_ca_w_2_400_s_0_360=1.01e-05
.param mcm4p1_cc_w_2_400_s_0_360=1.27e-10
.param mcm4p1_cf_w_2_400_s_0_360=1.84e-12
.param mcm4p1_ca_w_2_400_s_0_450=1.01e-05
.param mcm4p1_cc_w_2_400_s_0_450=1.15e-10
.param mcm4p1_cf_w_2_400_s_0_450=2.28e-12
.param mcm4p1_ca_w_2_400_s_0_600=1.01e-05
.param mcm4p1_cc_w_2_400_s_0_600=1.01e-10
.param mcm4p1_cf_w_2_400_s_0_600=3.01e-12
.param mcm4p1_ca_w_2_400_s_0_800=1.01e-05
.param mcm4p1_cc_w_2_400_s_0_800=8.61e-11
.param mcm4p1_cf_w_2_400_s_0_800=3.96e-12
.param mcm4p1_ca_w_2_400_s_1_000=1.01e-05
.param mcm4p1_cc_w_2_400_s_1_000=7.52e-11
.param mcm4p1_cf_w_2_400_s_1_000=4.89e-12
.param mcm4p1_ca_w_2_400_s_1_200=1.01e-05
.param mcm4p1_cc_w_2_400_s_1_200=6.70e-11
.param mcm4p1_cf_w_2_400_s_1_200=5.81e-12
.param mcm4p1_ca_w_2_400_s_2_100=1.01e-05
.param mcm4p1_cc_w_2_400_s_2_100=4.61e-11
.param mcm4p1_cf_w_2_400_s_2_100=9.67e-12
.param mcm4p1_ca_w_2_400_s_3_300=1.01e-05
.param mcm4p1_cc_w_2_400_s_3_300=3.29e-11
.param mcm4p1_cf_w_2_400_s_3_300=1.42e-11
.param mcm4p1_ca_w_2_400_s_9_000=1.01e-05
.param mcm4p1_cc_w_2_400_s_9_000=1.17e-11
.param mcm4p1_cf_w_2_400_s_9_000=2.75e-11
.param mcm4l1_ca_w_0_300_s_0_300=1.17e-05
.param mcm4l1_cc_w_0_300_s_0_300=1.08e-10
.param mcm4l1_cf_w_0_300_s_0_300=1.73e-12
.param mcm4l1_ca_w_0_300_s_0_360=1.17e-05
.param mcm4l1_cc_w_0_300_s_0_360=1.00e-10
.param mcm4l1_cf_w_0_300_s_0_360=2.07e-12
.param mcm4l1_ca_w_0_300_s_0_450=1.17e-05
.param mcm4l1_cc_w_0_300_s_0_450=9.07e-11
.param mcm4l1_cf_w_0_300_s_0_450=2.60e-12
.param mcm4l1_ca_w_0_300_s_0_600=1.17e-05
.param mcm4l1_cc_w_0_300_s_0_600=7.85e-11
.param mcm4l1_cf_w_0_300_s_0_600=3.46e-12
.param mcm4l1_ca_w_0_300_s_0_800=1.17e-05
.param mcm4l1_cc_w_0_300_s_0_800=6.65e-11
.param mcm4l1_cf_w_0_300_s_0_800=4.48e-12
.param mcm4l1_ca_w_0_300_s_1_000=1.17e-05
.param mcm4l1_cc_w_0_300_s_1_000=5.76e-11
.param mcm4l1_cf_w_0_300_s_1_000=5.53e-12
.param mcm4l1_ca_w_0_300_s_1_200=1.17e-05
.param mcm4l1_cc_w_0_300_s_1_200=5.08e-11
.param mcm4l1_cf_w_0_300_s_1_200=6.55e-12
.param mcm4l1_ca_w_0_300_s_2_100=1.17e-05
.param mcm4l1_cc_w_0_300_s_2_100=3.38e-11
.param mcm4l1_cf_w_0_300_s_2_100=1.10e-11
.param mcm4l1_ca_w_0_300_s_3_300=1.17e-05
.param mcm4l1_cc_w_0_300_s_3_300=2.35e-11
.param mcm4l1_cf_w_0_300_s_3_300=1.55e-11
.param mcm4l1_ca_w_0_300_s_9_000=1.17e-05
.param mcm4l1_cc_w_0_300_s_9_000=7.13e-12
.param mcm4l1_cf_w_0_300_s_9_000=2.73e-11
.param mcm4l1_ca_w_2_400_s_0_300=1.17e-05
.param mcm4l1_cc_w_2_400_s_0_300=1.34e-10
.param mcm4l1_cf_w_2_400_s_0_300=1.75e-12
.param mcm4l1_ca_w_2_400_s_0_360=1.17e-05
.param mcm4l1_cc_w_2_400_s_0_360=1.25e-10
.param mcm4l1_cf_w_2_400_s_0_360=2.09e-12
.param mcm4l1_ca_w_2_400_s_0_450=1.17e-05
.param mcm4l1_cc_w_2_400_s_0_450=1.14e-10
.param mcm4l1_cf_w_2_400_s_0_450=2.60e-12
.param mcm4l1_ca_w_2_400_s_0_600=1.17e-05
.param mcm4l1_cc_w_2_400_s_0_600=9.95e-11
.param mcm4l1_cf_w_2_400_s_0_600=3.43e-12
.param mcm4l1_ca_w_2_400_s_0_800=1.17e-05
.param mcm4l1_cc_w_2_400_s_0_800=8.47e-11
.param mcm4l1_cf_w_2_400_s_0_800=4.52e-12
.param mcm4l1_ca_w_2_400_s_1_000=1.17e-05
.param mcm4l1_cc_w_2_400_s_1_000=7.38e-11
.param mcm4l1_cf_w_2_400_s_1_000=5.58e-12
.param mcm4l1_ca_w_2_400_s_1_200=1.17e-05
.param mcm4l1_cc_w_2_400_s_1_200=6.56e-11
.param mcm4l1_cf_w_2_400_s_1_200=6.62e-12
.param mcm4l1_ca_w_2_400_s_2_100=1.17e-05
.param mcm4l1_cc_w_2_400_s_2_100=4.47e-11
.param mcm4l1_cf_w_2_400_s_2_100=1.10e-11
.param mcm4l1_ca_w_2_400_s_3_300=1.17e-05
.param mcm4l1_cc_w_2_400_s_3_300=3.14e-11
.param mcm4l1_cf_w_2_400_s_3_300=1.60e-11
.param mcm4l1_ca_w_2_400_s_9_000=1.17e-05
.param mcm4l1_cc_w_2_400_s_9_000=1.07e-11
.param mcm4l1_cf_w_2_400_s_9_000=2.98e-11
.param mcm4m1_ca_w_0_300_s_0_300=1.51e-05
.param mcm4m1_cc_w_0_300_s_0_300=1.06e-10
.param mcm4m1_cf_w_0_300_s_0_300=2.22e-12
.param mcm4m1_ca_w_0_300_s_0_360=1.51e-05
.param mcm4m1_cc_w_0_300_s_0_360=9.94e-11
.param mcm4m1_cf_w_0_300_s_0_360=2.65e-12
.param mcm4m1_ca_w_0_300_s_0_450=1.51e-05
.param mcm4m1_cc_w_0_300_s_0_450=8.98e-11
.param mcm4m1_cf_w_0_300_s_0_450=3.32e-12
.param mcm4m1_ca_w_0_300_s_0_600=1.51e-05
.param mcm4m1_cc_w_0_300_s_0_600=7.73e-11
.param mcm4m1_cf_w_0_300_s_0_600=4.40e-12
.param mcm4m1_ca_w_0_300_s_0_800=1.51e-05
.param mcm4m1_cc_w_0_300_s_0_800=6.51e-11
.param mcm4m1_cf_w_0_300_s_0_800=5.70e-12
.param mcm4m1_ca_w_0_300_s_1_000=1.51e-05
.param mcm4m1_cc_w_0_300_s_1_000=5.61e-11
.param mcm4m1_cf_w_0_300_s_1_000=7.02e-12
.param mcm4m1_ca_w_0_300_s_1_200=1.51e-05
.param mcm4m1_cc_w_0_300_s_1_200=4.92e-11
.param mcm4m1_cf_w_0_300_s_1_200=8.29e-12
.param mcm4m1_ca_w_0_300_s_2_100=1.51e-05
.param mcm4m1_cc_w_0_300_s_2_100=3.18e-11
.param mcm4m1_cf_w_0_300_s_2_100=1.37e-11
.param mcm4m1_ca_w_0_300_s_3_300=1.51e-05
.param mcm4m1_cc_w_0_300_s_3_300=2.14e-11
.param mcm4m1_cf_w_0_300_s_3_300=1.89e-11
.param mcm4m1_ca_w_0_300_s_9_000=1.51e-05
.param mcm4m1_cc_w_0_300_s_9_000=5.86e-12
.param mcm4m1_cf_w_0_300_s_9_000=3.09e-11
.param mcm4m1_ca_w_2_400_s_0_300=1.51e-05
.param mcm4m1_cc_w_2_400_s_0_300=1.32e-10
.param mcm4m1_cf_w_2_400_s_0_300=2.23e-12
.param mcm4m1_ca_w_2_400_s_0_360=1.51e-05
.param mcm4m1_cc_w_2_400_s_0_360=1.23e-10
.param mcm4m1_cf_w_2_400_s_0_360=2.66e-12
.param mcm4m1_ca_w_2_400_s_0_450=1.51e-05
.param mcm4m1_cc_w_2_400_s_0_450=1.12e-10
.param mcm4m1_cf_w_2_400_s_0_450=3.31e-12
.param mcm4m1_ca_w_2_400_s_0_600=1.51e-05
.param mcm4m1_cc_w_2_400_s_0_600=9.70e-11
.param mcm4m1_cf_w_2_400_s_0_600=4.36e-12
.param mcm4m1_ca_w_2_400_s_0_800=1.51e-05
.param mcm4m1_cc_w_2_400_s_0_800=8.21e-11
.param mcm4m1_cf_w_2_400_s_0_800=5.74e-12
.param mcm4m1_ca_w_2_400_s_1_000=1.51e-05
.param mcm4m1_cc_w_2_400_s_1_000=7.12e-11
.param mcm4m1_cf_w_2_400_s_1_000=7.07e-12
.param mcm4m1_ca_w_2_400_s_1_200=1.51e-05
.param mcm4m1_cc_w_2_400_s_1_200=6.30e-11
.param mcm4m1_cf_w_2_400_s_1_200=8.35e-12
.param mcm4m1_ca_w_2_400_s_2_100=1.51e-05
.param mcm4m1_cc_w_2_400_s_2_100=4.21e-11
.param mcm4m1_cf_w_2_400_s_2_100=1.36e-11
.param mcm4m1_ca_w_2_400_s_3_300=1.51e-05
.param mcm4m1_cc_w_2_400_s_3_300=2.89e-11
.param mcm4m1_cf_w_2_400_s_3_300=1.95e-11
.param mcm4m1_ca_w_2_400_s_9_000=1.51e-05
.param mcm4m1_cc_w_2_400_s_9_000=9.10e-12
.param mcm4m1_cf_w_2_400_s_9_000=3.39e-11
.param mcm4m2_ca_w_0_300_s_0_300=2.09e-05
.param mcm4m2_cc_w_0_300_s_0_300=1.05e-10
.param mcm4m2_cf_w_0_300_s_0_300=3.04e-12
.param mcm4m2_ca_w_0_300_s_0_360=2.09e-05
.param mcm4m2_cc_w_0_300_s_0_360=9.77e-11
.param mcm4m2_cf_w_0_300_s_0_360=3.63e-12
.param mcm4m2_ca_w_0_300_s_0_450=2.09e-05
.param mcm4m2_cc_w_0_300_s_0_450=8.80e-11
.param mcm4m2_cf_w_0_300_s_0_450=4.52e-12
.param mcm4m2_ca_w_0_300_s_0_600=2.09e-05
.param mcm4m2_cc_w_0_300_s_0_600=7.54e-11
.param mcm4m2_cf_w_0_300_s_0_600=5.97e-12
.param mcm4m2_ca_w_0_300_s_0_800=2.09e-05
.param mcm4m2_cc_w_0_300_s_0_800=6.31e-11
.param mcm4m2_cf_w_0_300_s_0_800=7.72e-12
.param mcm4m2_ca_w_0_300_s_1_000=2.09e-05
.param mcm4m2_cc_w_0_300_s_1_000=5.38e-11
.param mcm4m2_cf_w_0_300_s_1_000=9.44e-12
.param mcm4m2_ca_w_0_300_s_1_200=2.09e-05
.param mcm4m2_cc_w_0_300_s_1_200=4.68e-11
.param mcm4m2_cf_w_0_300_s_1_200=1.11e-11
.param mcm4m2_ca_w_0_300_s_2_100=2.09e-05
.param mcm4m2_cc_w_0_300_s_2_100=2.90e-11
.param mcm4m2_cf_w_0_300_s_2_100=1.78e-11
.param mcm4m2_ca_w_0_300_s_3_300=2.09e-05
.param mcm4m2_cc_w_0_300_s_3_300=1.88e-11
.param mcm4m2_cf_w_0_300_s_3_300=2.38e-11
.param mcm4m2_ca_w_0_300_s_9_000=2.09e-05
.param mcm4m2_cc_w_0_300_s_9_000=4.49e-12
.param mcm4m2_cf_w_0_300_s_9_000=3.56e-11
.param mcm4m2_ca_w_2_400_s_0_300=2.09e-05
.param mcm4m2_cc_w_2_400_s_0_300=1.28e-10
.param mcm4m2_cf_w_2_400_s_0_300=3.05e-12
.param mcm4m2_ca_w_2_400_s_0_360=2.09e-05
.param mcm4m2_cc_w_2_400_s_0_360=1.20e-10
.param mcm4m2_cf_w_2_400_s_0_360=3.64e-12
.param mcm4m2_ca_w_2_400_s_0_450=2.09e-05
.param mcm4m2_cc_w_2_400_s_0_450=1.08e-10
.param mcm4m2_cf_w_2_400_s_0_450=4.52e-12
.param mcm4m2_ca_w_2_400_s_0_600=2.09e-05
.param mcm4m2_cc_w_2_400_s_0_600=9.36e-11
.param mcm4m2_cf_w_2_400_s_0_600=5.93e-12
.param mcm4m2_ca_w_2_400_s_0_800=2.09e-05
.param mcm4m2_cc_w_2_400_s_0_800=7.88e-11
.param mcm4m2_cf_w_2_400_s_0_800=7.76e-12
.param mcm4m2_ca_w_2_400_s_1_000=2.09e-05
.param mcm4m2_cc_w_2_400_s_1_000=6.78e-11
.param mcm4m2_cf_w_2_400_s_1_000=9.53e-12
.param mcm4m2_ca_w_2_400_s_1_200=2.09e-05
.param mcm4m2_cc_w_2_400_s_1_200=5.95e-11
.param mcm4m2_cf_w_2_400_s_1_200=1.12e-11
.param mcm4m2_ca_w_2_400_s_2_100=2.09e-05
.param mcm4m2_cc_w_2_400_s_2_100=3.89e-11
.param mcm4m2_cf_w_2_400_s_2_100=1.78e-11
.param mcm4m2_ca_w_2_400_s_3_300=2.09e-05
.param mcm4m2_cc_w_2_400_s_3_300=2.59e-11
.param mcm4m2_cf_w_2_400_s_3_300=2.46e-11
.param mcm4m2_ca_w_2_400_s_9_000=2.09e-05
.param mcm4m2_cc_w_2_400_s_9_000=7.40e-12
.param mcm4m2_cf_w_2_400_s_9_000=3.92e-11
.param mcm4m3_ca_w_0_300_s_0_300=8.85e-05
.param mcm4m3_cc_w_0_300_s_0_300=9.36e-11
.param mcm4m3_cf_w_0_300_s_0_300=1.18e-11
.param mcm4m3_ca_w_0_300_s_0_360=8.85e-05
.param mcm4m3_cc_w_0_300_s_0_360=8.61e-11
.param mcm4m3_cf_w_0_300_s_0_360=1.39e-11
.param mcm4m3_ca_w_0_300_s_0_450=8.85e-05
.param mcm4m3_cc_w_0_300_s_0_450=7.62e-11
.param mcm4m3_cf_w_0_300_s_0_450=1.67e-11
.param mcm4m3_ca_w_0_300_s_0_600=8.85e-05
.param mcm4m3_cc_w_0_300_s_0_600=6.30e-11
.param mcm4m3_cf_w_0_300_s_0_600=2.11e-11
.param mcm4m3_ca_w_0_300_s_0_800=8.85e-05
.param mcm4m3_cc_w_0_300_s_0_800=5.05e-11
.param mcm4m3_cf_w_0_300_s_0_800=2.58e-11
.param mcm4m3_ca_w_0_300_s_1_000=8.85e-05
.param mcm4m3_cc_w_0_300_s_1_000=4.13e-11
.param mcm4m3_cf_w_0_300_s_1_000=2.99e-11
.param mcm4m3_ca_w_0_300_s_1_200=8.85e-05
.param mcm4m3_cc_w_0_300_s_1_200=3.45e-11
.param mcm4m3_cf_w_0_300_s_1_200=3.34e-11
.param mcm4m3_ca_w_0_300_s_2_100=8.85e-05
.param mcm4m3_cc_w_0_300_s_2_100=1.80e-11
.param mcm4m3_cf_w_0_300_s_2_100=4.46e-11
.param mcm4m3_ca_w_0_300_s_3_300=8.85e-05
.param mcm4m3_cc_w_0_300_s_3_300=1.01e-11
.param mcm4m3_cf_w_0_300_s_3_300=5.12e-11
.param mcm4m3_ca_w_0_300_s_9_000=8.85e-05
.param mcm4m3_cc_w_0_300_s_9_000=1.90e-12
.param mcm4m3_cf_w_0_300_s_9_000=5.91e-11
.param mcm4m3_ca_w_2_400_s_0_300=8.85e-05
.param mcm4m3_cc_w_2_400_s_0_300=1.12e-10
.param mcm4m3_cf_w_2_400_s_0_300=1.18e-11
.param mcm4m3_ca_w_2_400_s_0_360=8.85e-05
.param mcm4m3_cc_w_2_400_s_0_360=1.04e-10
.param mcm4m3_cf_w_2_400_s_0_360=1.39e-11
.param mcm4m3_ca_w_2_400_s_0_450=8.85e-05
.param mcm4m3_cc_w_2_400_s_0_450=9.29e-11
.param mcm4m3_cf_w_2_400_s_0_450=1.68e-11
.param mcm4m3_ca_w_2_400_s_0_600=8.85e-05
.param mcm4m3_cc_w_2_400_s_0_600=7.84e-11
.param mcm4m3_cf_w_2_400_s_0_600=2.10e-11
.param mcm4m3_ca_w_2_400_s_0_800=8.85e-05
.param mcm4m3_cc_w_2_400_s_0_800=6.42e-11
.param mcm4m3_cf_w_2_400_s_0_800=2.59e-11
.param mcm4m3_ca_w_2_400_s_1_000=8.85e-05
.param mcm4m3_cc_w_2_400_s_1_000=5.38e-11
.param mcm4m3_cf_w_2_400_s_1_000=3.00e-11
.param mcm4m3_ca_w_2_400_s_1_200=8.85e-05
.param mcm4m3_cc_w_2_400_s_1_200=4.61e-11
.param mcm4m3_cf_w_2_400_s_1_200=3.35e-11
.param mcm4m3_ca_w_2_400_s_2_100=8.85e-05
.param mcm4m3_cc_w_2_400_s_2_100=2.75e-11
.param mcm4m3_cf_w_2_400_s_2_100=4.46e-11
.param mcm4m3_ca_w_2_400_s_3_300=8.85e-05
.param mcm4m3_cc_w_2_400_s_3_300=1.67e-11
.param mcm4m3_cf_w_2_400_s_3_300=5.31e-11
.param mcm4m3_ca_w_2_400_s_9_000=8.85e-05
.param mcm4m3_cc_w_2_400_s_9_000=3.95e-12
.param mcm4m3_cf_w_2_400_s_9_000=6.50e-11
.param mcm5f_ca_w_1_600_s_1_600=6.48e-06
.param mcm5f_cc_w_1_600_s_1_600=7.35e-11
.param mcm5f_cf_w_1_600_s_1_600=5.01e-12
.param mcm5f_ca_w_1_600_s_1_700=6.48e-06
.param mcm5f_cc_w_1_600_s_1_700=6.99e-11
.param mcm5f_cf_w_1_600_s_1_700=5.31e-12
.param mcm5f_ca_w_1_600_s_1_900=6.48e-06
.param mcm5f_cc_w_1_600_s_1_900=6.37e-11
.param mcm5f_cf_w_1_600_s_1_900=5.90e-12
.param mcm5f_ca_w_1_600_s_2_000=6.48e-06
.param mcm5f_cc_w_1_600_s_2_000=6.11e-11
.param mcm5f_cf_w_1_600_s_2_000=6.19e-12
.param mcm5f_ca_w_1_600_s_2_400=6.48e-06
.param mcm5f_cc_w_1_600_s_2_400=5.27e-11
.param mcm5f_cf_w_1_600_s_2_400=7.34e-12
.param mcm5f_ca_w_1_600_s_2_800=6.48e-06
.param mcm5f_cc_w_1_600_s_2_800=4.65e-11
.param mcm5f_cf_w_1_600_s_2_800=8.47e-12
.param mcm5f_ca_w_1_600_s_3_200=6.48e-06
.param mcm5f_cc_w_1_600_s_3_200=4.18e-11
.param mcm5f_cf_w_1_600_s_3_200=9.54e-12
.param mcm5f_ca_w_1_600_s_4_800=6.48e-06
.param mcm5f_cc_w_1_600_s_4_800=2.97e-11
.param mcm5f_cf_w_1_600_s_4_800=1.35e-11
.param mcm5f_ca_w_1_600_s_10_000=6.48e-06
.param mcm5f_cc_w_1_600_s_10_000=1.40e-11
.param mcm5f_cf_w_1_600_s_10_000=2.27e-11
.param mcm5f_ca_w_1_600_s_12_000=6.48e-06
.param mcm5f_cc_w_1_600_s_12_000=1.11e-11
.param mcm5f_cf_w_1_600_s_12_000=2.50e-11
.param mcm5f_ca_w_4_000_s_1_600=6.48e-06
.param mcm5f_cc_w_4_000_s_1_600=8.04e-11
.param mcm5f_cf_w_4_000_s_1_600=5.02e-12
.param mcm5f_ca_w_4_000_s_1_700=6.48e-06
.param mcm5f_cc_w_4_000_s_1_700=7.64e-11
.param mcm5f_cf_w_4_000_s_1_700=5.32e-12
.param mcm5f_ca_w_4_000_s_1_900=6.48e-06
.param mcm5f_cc_w_4_000_s_1_900=6.99e-11
.param mcm5f_cf_w_4_000_s_1_900=5.91e-12
.param mcm5f_ca_w_4_000_s_2_000=6.48e-06
.param mcm5f_cc_w_4_000_s_2_000=6.72e-11
.param mcm5f_cf_w_4_000_s_2_000=6.20e-12
.param mcm5f_ca_w_4_000_s_2_400=6.48e-06
.param mcm5f_cc_w_4_000_s_2_400=5.83e-11
.param mcm5f_cf_w_4_000_s_2_400=7.35e-12
.param mcm5f_ca_w_4_000_s_2_800=6.48e-06
.param mcm5f_cc_w_4_000_s_2_800=5.18e-11
.param mcm5f_cf_w_4_000_s_2_800=8.48e-12
.param mcm5f_ca_w_4_000_s_3_200=6.48e-06
.param mcm5f_cc_w_4_000_s_3_200=4.67e-11
.param mcm5f_cf_w_4_000_s_3_200=9.57e-12
.param mcm5f_ca_w_4_000_s_4_800=6.48e-06
.param mcm5f_cc_w_4_000_s_4_800=3.36e-11
.param mcm5f_cf_w_4_000_s_4_800=1.36e-11
.param mcm5f_ca_w_4_000_s_10_000=6.48e-06
.param mcm5f_cc_w_4_000_s_10_000=1.66e-11
.param mcm5f_cf_w_4_000_s_10_000=2.31e-11
.param mcm5f_ca_w_4_000_s_12_000=6.48e-06
.param mcm5f_cc_w_4_000_s_12_000=1.34e-11
.param mcm5f_cf_w_4_000_s_12_000=2.56e-11
.param mcm5d_ca_w_1_600_s_1_600=6.88e-06
.param mcm5d_cc_w_1_600_s_1_600=7.31e-11
.param mcm5d_cf_w_1_600_s_1_600=5.31e-12
.param mcm5d_ca_w_1_600_s_1_700=6.88e-06
.param mcm5d_cc_w_1_600_s_1_700=6.95e-11
.param mcm5d_cf_w_1_600_s_1_700=5.62e-12
.param mcm5d_ca_w_1_600_s_1_900=6.88e-06
.param mcm5d_cc_w_1_600_s_1_900=6.32e-11
.param mcm5d_cf_w_1_600_s_1_900=6.25e-12
.param mcm5d_ca_w_1_600_s_2_000=6.88e-06
.param mcm5d_cc_w_1_600_s_2_000=6.06e-11
.param mcm5d_cf_w_1_600_s_2_000=6.56e-12
.param mcm5d_ca_w_1_600_s_2_400=6.88e-06
.param mcm5d_cc_w_1_600_s_2_400=5.22e-11
.param mcm5d_cf_w_1_600_s_2_400=7.77e-12
.param mcm5d_ca_w_1_600_s_2_800=6.88e-06
.param mcm5d_cc_w_1_600_s_2_800=4.60e-11
.param mcm5d_cf_w_1_600_s_2_800=8.95e-12
.param mcm5d_ca_w_1_600_s_3_200=6.88e-06
.param mcm5d_cc_w_1_600_s_3_200=4.13e-11
.param mcm5d_cf_w_1_600_s_3_200=1.01e-11
.param mcm5d_ca_w_1_600_s_4_800=6.88e-06
.param mcm5d_cc_w_1_600_s_4_800=2.91e-11
.param mcm5d_cf_w_1_600_s_4_800=1.42e-11
.param mcm5d_ca_w_1_600_s_10_000=6.88e-06
.param mcm5d_cc_w_1_600_s_10_000=1.35e-11
.param mcm5d_cf_w_1_600_s_10_000=2.36e-11
.param mcm5d_ca_w_1_600_s_12_000=6.88e-06
.param mcm5d_cc_w_1_600_s_12_000=1.07e-11
.param mcm5d_cf_w_1_600_s_12_000=2.59e-11
.param mcm5d_ca_w_4_000_s_1_600=6.88e-06
.param mcm5d_cc_w_4_000_s_1_600=7.98e-11
.param mcm5d_cf_w_4_000_s_1_600=5.31e-12
.param mcm5d_ca_w_4_000_s_1_700=6.88e-06
.param mcm5d_cc_w_4_000_s_1_700=7.59e-11
.param mcm5d_cf_w_4_000_s_1_700=5.63e-12
.param mcm5d_ca_w_4_000_s_1_900=6.88e-06
.param mcm5d_cc_w_4_000_s_1_900=6.94e-11
.param mcm5d_cf_w_4_000_s_1_900=6.26e-12
.param mcm5d_ca_w_4_000_s_2_000=6.88e-06
.param mcm5d_cc_w_4_000_s_2_000=6.66e-11
.param mcm5d_cf_w_4_000_s_2_000=6.57e-12
.param mcm5d_ca_w_4_000_s_2_400=6.88e-06
.param mcm5d_cc_w_4_000_s_2_400=5.77e-11
.param mcm5d_cf_w_4_000_s_2_400=7.78e-12
.param mcm5d_ca_w_4_000_s_2_800=6.88e-06
.param mcm5d_cc_w_4_000_s_2_800=5.12e-11
.param mcm5d_cf_w_4_000_s_2_800=8.97e-12
.param mcm5d_ca_w_4_000_s_3_200=6.88e-06
.param mcm5d_cc_w_4_000_s_3_200=4.61e-11
.param mcm5d_cf_w_4_000_s_3_200=1.01e-11
.param mcm5d_ca_w_4_000_s_4_800=6.88e-06
.param mcm5d_cc_w_4_000_s_4_800=3.30e-11
.param mcm5d_cf_w_4_000_s_4_800=1.43e-11
.param mcm5d_ca_w_4_000_s_10_000=6.88e-06
.param mcm5d_cc_w_4_000_s_10_000=1.61e-11
.param mcm5d_cf_w_4_000_s_10_000=2.41e-11
.param mcm5d_ca_w_4_000_s_12_000=6.88e-06
.param mcm5d_cc_w_4_000_s_12_000=1.30e-11
.param mcm5d_cf_w_4_000_s_12_000=2.65e-11
.param mcm5p1_ca_w_1_600_s_1_600=7.26e-06
.param mcm5p1_cc_w_1_600_s_1_600=7.27e-11
.param mcm5p1_cf_w_1_600_s_1_600=5.59e-12
.param mcm5p1_ca_w_1_600_s_1_700=7.26e-06
.param mcm5p1_cc_w_1_600_s_1_700=6.91e-11
.param mcm5p1_cf_w_1_600_s_1_700=5.92e-12
.param mcm5p1_ca_w_1_600_s_1_900=7.26e-06
.param mcm5p1_cc_w_1_600_s_1_900=6.28e-11
.param mcm5p1_cf_w_1_600_s_1_900=6.58e-12
.param mcm5p1_ca_w_1_600_s_2_000=7.26e-06
.param mcm5p1_cc_w_1_600_s_2_000=6.02e-11
.param mcm5p1_cf_w_1_600_s_2_000=6.91e-12
.param mcm5p1_ca_w_1_600_s_2_400=7.26e-06
.param mcm5p1_cc_w_1_600_s_2_400=5.18e-11
.param mcm5p1_cf_w_1_600_s_2_400=8.18e-12
.param mcm5p1_ca_w_1_600_s_2_800=7.26e-06
.param mcm5p1_cc_w_1_600_s_2_800=4.56e-11
.param mcm5p1_cf_w_1_600_s_2_800=9.41e-12
.param mcm5p1_ca_w_1_600_s_3_200=7.26e-06
.param mcm5p1_cc_w_1_600_s_3_200=4.08e-11
.param mcm5p1_cf_w_1_600_s_3_200=1.06e-11
.param mcm5p1_ca_w_1_600_s_4_800=7.26e-06
.param mcm5p1_cc_w_1_600_s_4_800=2.86e-11
.param mcm5p1_cf_w_1_600_s_4_800=1.49e-11
.param mcm5p1_ca_w_1_600_s_10_000=7.26e-06
.param mcm5p1_cc_w_1_600_s_10_000=1.31e-11
.param mcm5p1_cf_w_1_600_s_10_000=2.45e-11
.param mcm5p1_ca_w_1_600_s_12_000=7.26e-06
.param mcm5p1_cc_w_1_600_s_12_000=1.03e-11
.param mcm5p1_cf_w_1_600_s_12_000=2.68e-11
.param mcm5p1_ca_w_4_000_s_1_600=7.26e-06
.param mcm5p1_cc_w_4_000_s_1_600=7.93e-11
.param mcm5p1_cf_w_4_000_s_1_600=5.61e-12
.param mcm5p1_ca_w_4_000_s_1_700=7.26e-06
.param mcm5p1_cc_w_4_000_s_1_700=7.54e-11
.param mcm5p1_cf_w_4_000_s_1_700=5.94e-12
.param mcm5p1_ca_w_4_000_s_1_900=7.26e-06
.param mcm5p1_cc_w_4_000_s_1_900=6.89e-11
.param mcm5p1_cf_w_4_000_s_1_900=6.59e-12
.param mcm5p1_ca_w_4_000_s_2_000=7.26e-06
.param mcm5p1_cc_w_4_000_s_2_000=6.62e-11
.param mcm5p1_cf_w_4_000_s_2_000=6.92e-12
.param mcm5p1_ca_w_4_000_s_2_400=7.26e-06
.param mcm5p1_cc_w_4_000_s_2_400=5.71e-11
.param mcm5p1_cf_w_4_000_s_2_400=8.19e-12
.param mcm5p1_ca_w_4_000_s_2_800=7.26e-06
.param mcm5p1_cc_w_4_000_s_2_800=5.06e-11
.param mcm5p1_cf_w_4_000_s_2_800=9.43e-12
.param mcm5p1_ca_w_4_000_s_3_200=7.26e-06
.param mcm5p1_cc_w_4_000_s_3_200=4.55e-11
.param mcm5p1_cf_w_4_000_s_3_200=1.06e-11
.param mcm5p1_ca_w_4_000_s_4_800=7.26e-06
.param mcm5p1_cc_w_4_000_s_4_800=3.25e-11
.param mcm5p1_cf_w_4_000_s_4_800=1.50e-11
.param mcm5p1_ca_w_4_000_s_10_000=7.26e-06
.param mcm5p1_cc_w_4_000_s_10_000=1.56e-11
.param mcm5p1_cf_w_4_000_s_10_000=2.49e-11
.param mcm5p1_ca_w_4_000_s_12_000=7.26e-06
.param mcm5p1_cc_w_4_000_s_12_000=1.26e-11
.param mcm5p1_cf_w_4_000_s_12_000=2.74e-11
.param mcm5l1_ca_w_1_600_s_1_600=8.04e-06
.param mcm5l1_cc_w_1_600_s_1_600=7.19e-11
.param mcm5l1_cf_w_1_600_s_1_600=6.16e-12
.param mcm5l1_ca_w_1_600_s_1_700=8.04e-06
.param mcm5l1_cc_w_1_600_s_1_700=6.82e-11
.param mcm5l1_cf_w_1_600_s_1_700=6.52e-12
.param mcm5l1_ca_w_1_600_s_1_900=8.04e-06
.param mcm5l1_cc_w_1_600_s_1_900=6.20e-11
.param mcm5l1_cf_w_1_600_s_1_900=7.24e-12
.param mcm5l1_ca_w_1_600_s_2_000=8.04e-06
.param mcm5l1_cc_w_1_600_s_2_000=5.94e-11
.param mcm5l1_cf_w_1_600_s_2_000=7.59e-12
.param mcm5l1_ca_w_1_600_s_2_400=8.04e-06
.param mcm5l1_cc_w_1_600_s_2_400=5.09e-11
.param mcm5l1_cf_w_1_600_s_2_400=8.98e-12
.param mcm5l1_ca_w_1_600_s_2_800=8.04e-06
.param mcm5l1_cc_w_1_600_s_2_800=4.47e-11
.param mcm5l1_cf_w_1_600_s_2_800=1.03e-11
.param mcm5l1_ca_w_1_600_s_3_200=8.04e-06
.param mcm5l1_cc_w_1_600_s_3_200=3.99e-11
.param mcm5l1_cf_w_1_600_s_3_200=1.16e-11
.param mcm5l1_ca_w_1_600_s_4_800=8.04e-06
.param mcm5l1_cc_w_1_600_s_4_800=2.77e-11
.param mcm5l1_cf_w_1_600_s_4_800=1.62e-11
.param mcm5l1_ca_w_1_600_s_10_000=8.04e-06
.param mcm5l1_cc_w_1_600_s_10_000=1.23e-11
.param mcm5l1_cf_w_1_600_s_10_000=2.61e-11
.param mcm5l1_ca_w_1_600_s_12_000=8.04e-06
.param mcm5l1_cc_w_1_600_s_12_000=9.59e-12
.param mcm5l1_cf_w_1_600_s_12_000=2.84e-11
.param mcm5l1_ca_w_4_000_s_1_600=8.04e-06
.param mcm5l1_cc_w_4_000_s_1_600=7.83e-11
.param mcm5l1_cf_w_4_000_s_1_600=6.16e-12
.param mcm5l1_ca_w_4_000_s_1_700=8.04e-06
.param mcm5l1_cc_w_4_000_s_1_700=7.44e-11
.param mcm5l1_cf_w_4_000_s_1_700=6.53e-12
.param mcm5l1_ca_w_4_000_s_1_900=8.04e-06
.param mcm5l1_cc_w_4_000_s_1_900=6.78e-11
.param mcm5l1_cf_w_4_000_s_1_900=7.25e-12
.param mcm5l1_ca_w_4_000_s_2_000=8.04e-06
.param mcm5l1_cc_w_4_000_s_2_000=6.51e-11
.param mcm5l1_cf_w_4_000_s_2_000=7.60e-12
.param mcm5l1_ca_w_4_000_s_2_400=8.04e-06
.param mcm5l1_cc_w_4_000_s_2_400=5.62e-11
.param mcm5l1_cf_w_4_000_s_2_400=9.00e-12
.param mcm5l1_ca_w_4_000_s_2_800=8.04e-06
.param mcm5l1_cc_w_4_000_s_2_800=4.96e-11
.param mcm5l1_cf_w_4_000_s_2_800=1.03e-11
.param mcm5l1_ca_w_4_000_s_3_200=8.04e-06
.param mcm5l1_cc_w_4_000_s_3_200=4.44e-11
.param mcm5l1_cf_w_4_000_s_3_200=1.16e-11
.param mcm5l1_ca_w_4_000_s_4_800=8.04e-06
.param mcm5l1_cc_w_4_000_s_4_800=3.15e-11
.param mcm5l1_cf_w_4_000_s_4_800=1.63e-11
.param mcm5l1_ca_w_4_000_s_10_000=8.04e-06
.param mcm5l1_cc_w_4_000_s_10_000=1.48e-11
.param mcm5l1_cf_w_4_000_s_10_000=2.66e-11
.param mcm5l1_ca_w_4_000_s_12_000=8.04e-06
.param mcm5l1_cc_w_4_000_s_12_000=1.18e-11
.param mcm5l1_cf_w_4_000_s_12_000=2.91e-11
.param mcm5m1_ca_w_1_600_s_1_600=9.50e-06
.param mcm5m1_cc_w_1_600_s_1_600=7.04e-11
.param mcm5m1_cf_w_1_600_s_1_600=7.21e-12
.param mcm5m1_ca_w_1_600_s_1_700=9.50e-06
.param mcm5m1_cc_w_1_600_s_1_700=6.68e-11
.param mcm5m1_cf_w_1_600_s_1_700=7.63e-12
.param mcm5m1_ca_w_1_600_s_1_900=9.50e-06
.param mcm5m1_cc_w_1_600_s_1_900=6.05e-11
.param mcm5m1_cf_w_1_600_s_1_900=8.47e-12
.param mcm5m1_ca_w_1_600_s_2_000=9.50e-06
.param mcm5m1_cc_w_1_600_s_2_000=5.79e-11
.param mcm5m1_cf_w_1_600_s_2_000=8.88e-12
.param mcm5m1_ca_w_1_600_s_2_400=9.50e-06
.param mcm5m1_cc_w_1_600_s_2_400=4.94e-11
.param mcm5m1_cf_w_1_600_s_2_400=1.05e-11
.param mcm5m1_ca_w_1_600_s_2_800=9.50e-06
.param mcm5m1_cc_w_1_600_s_2_800=4.32e-11
.param mcm5m1_cf_w_1_600_s_2_800=1.20e-11
.param mcm5m1_ca_w_1_600_s_3_200=9.50e-06
.param mcm5m1_cc_w_1_600_s_3_200=3.84e-11
.param mcm5m1_cf_w_1_600_s_3_200=1.35e-11
.param mcm5m1_ca_w_1_600_s_4_800=9.50e-06
.param mcm5m1_cc_w_1_600_s_4_800=2.61e-11
.param mcm5m1_cf_w_1_600_s_4_800=1.86e-11
.param mcm5m1_ca_w_1_600_s_10_000=9.50e-06
.param mcm5m1_cc_w_1_600_s_10_000=1.10e-11
.param mcm5m1_cf_w_1_600_s_10_000=2.90e-11
.param mcm5m1_ca_w_1_600_s_12_000=9.50e-06
.param mcm5m1_cc_w_1_600_s_12_000=8.51e-12
.param mcm5m1_cf_w_1_600_s_12_000=3.11e-11
.param mcm5m1_ca_w_4_000_s_1_600=9.50e-06
.param mcm5m1_cc_w_4_000_s_1_600=7.66e-11
.param mcm5m1_cf_w_4_000_s_1_600=7.22e-12
.param mcm5m1_ca_w_4_000_s_1_700=9.50e-06
.param mcm5m1_cc_w_4_000_s_1_700=7.27e-11
.param mcm5m1_cf_w_4_000_s_1_700=7.64e-12
.param mcm5m1_ca_w_4_000_s_1_900=9.50e-06
.param mcm5m1_cc_w_4_000_s_1_900=6.61e-11
.param mcm5m1_cf_w_4_000_s_1_900=8.47e-12
.param mcm5m1_ca_w_4_000_s_2_000=9.50e-06
.param mcm5m1_cc_w_4_000_s_2_000=6.33e-11
.param mcm5m1_cf_w_4_000_s_2_000=8.88e-12
.param mcm5m1_ca_w_4_000_s_2_400=9.50e-06
.param mcm5m1_cc_w_4_000_s_2_400=5.45e-11
.param mcm5m1_cf_w_4_000_s_2_400=1.05e-11
.param mcm5m1_ca_w_4_000_s_2_800=9.50e-06
.param mcm5m1_cc_w_4_000_s_2_800=4.78e-11
.param mcm5m1_cf_w_4_000_s_2_800=1.20e-11
.param mcm5m1_ca_w_4_000_s_3_200=9.50e-06
.param mcm5m1_cc_w_4_000_s_3_200=4.27e-11
.param mcm5m1_cf_w_4_000_s_3_200=1.35e-11
.param mcm5m1_ca_w_4_000_s_4_800=9.50e-06
.param mcm5m1_cc_w_4_000_s_4_800=2.98e-11
.param mcm5m1_cf_w_4_000_s_4_800=1.87e-11
.param mcm5m1_ca_w_4_000_s_10_000=9.50e-06
.param mcm5m1_cc_w_4_000_s_10_000=1.35e-11
.param mcm5m1_cf_w_4_000_s_10_000=2.95e-11
.param mcm5m1_ca_w_4_000_s_12_000=9.50e-06
.param mcm5m1_cc_w_4_000_s_12_000=1.07e-11
.param mcm5m1_cf_w_4_000_s_12_000=3.19e-11
.param mcm5m2_ca_w_1_600_s_1_600=1.15e-05
.param mcm5m2_cc_w_1_600_s_1_600=6.87e-11
.param mcm5m2_cf_w_1_600_s_1_600=8.63e-12
.param mcm5m2_ca_w_1_600_s_1_700=1.15e-05
.param mcm5m2_cc_w_1_600_s_1_700=6.51e-11
.param mcm5m2_cf_w_1_600_s_1_700=9.13e-12
.param mcm5m2_ca_w_1_600_s_1_900=1.15e-05
.param mcm5m2_cc_w_1_600_s_1_900=5.88e-11
.param mcm5m2_cf_w_1_600_s_1_900=1.01e-11
.param mcm5m2_ca_w_1_600_s_2_000=1.15e-05
.param mcm5m2_cc_w_1_600_s_2_000=5.61e-11
.param mcm5m2_cf_w_1_600_s_2_000=1.06e-11
.param mcm5m2_ca_w_1_600_s_2_400=1.15e-05
.param mcm5m2_cc_w_1_600_s_2_400=4.77e-11
.param mcm5m2_cf_w_1_600_s_2_400=1.24e-11
.param mcm5m2_ca_w_1_600_s_2_800=1.15e-05
.param mcm5m2_cc_w_1_600_s_2_800=4.14e-11
.param mcm5m2_cf_w_1_600_s_2_800=1.42e-11
.param mcm5m2_ca_w_1_600_s_3_200=1.15e-05
.param mcm5m2_cc_w_1_600_s_3_200=3.65e-11
.param mcm5m2_cf_w_1_600_s_3_200=1.59e-11
.param mcm5m2_ca_w_1_600_s_4_800=1.15e-05
.param mcm5m2_cc_w_1_600_s_4_800=2.43e-11
.param mcm5m2_cf_w_1_600_s_4_800=2.16e-11
.param mcm5m2_ca_w_1_600_s_10_000=1.15e-05
.param mcm5m2_cc_w_1_600_s_10_000=9.75e-12
.param mcm5m2_cf_w_1_600_s_10_000=3.23e-11
.param mcm5m2_ca_w_1_600_s_12_000=1.15e-05
.param mcm5m2_cc_w_1_600_s_12_000=7.42e-12
.param mcm5m2_cf_w_1_600_s_12_000=3.44e-11
.param mcm5m2_ca_w_4_000_s_1_600=1.15e-05
.param mcm5m2_cc_w_4_000_s_1_600=7.45e-11
.param mcm5m2_cf_w_4_000_s_1_600=8.63e-12
.param mcm5m2_ca_w_4_000_s_1_700=1.15e-05
.param mcm5m2_cc_w_4_000_s_1_700=7.06e-11
.param mcm5m2_cf_w_4_000_s_1_700=9.13e-12
.param mcm5m2_ca_w_4_000_s_1_900=1.15e-05
.param mcm5m2_cc_w_4_000_s_1_900=6.41e-11
.param mcm5m2_cf_w_4_000_s_1_900=1.01e-11
.param mcm5m2_ca_w_4_000_s_2_000=1.15e-05
.param mcm5m2_cc_w_4_000_s_2_000=6.13e-11
.param mcm5m2_cf_w_4_000_s_2_000=1.06e-11
.param mcm5m2_ca_w_4_000_s_2_400=1.15e-05
.param mcm5m2_cc_w_4_000_s_2_400=5.25e-11
.param mcm5m2_cf_w_4_000_s_2_400=1.25e-11
.param mcm5m2_ca_w_4_000_s_2_800=1.15e-05
.param mcm5m2_cc_w_4_000_s_2_800=4.59e-11
.param mcm5m2_cf_w_4_000_s_2_800=1.42e-11
.param mcm5m2_ca_w_4_000_s_3_200=1.15e-05
.param mcm5m2_cc_w_4_000_s_3_200=4.07e-11
.param mcm5m2_cf_w_4_000_s_3_200=1.59e-11
.param mcm5m2_ca_w_4_000_s_4_800=1.15e-05
.param mcm5m2_cc_w_4_000_s_4_800=2.79e-11
.param mcm5m2_cf_w_4_000_s_4_800=2.17e-11
.param mcm5m2_ca_w_4_000_s_10_000=1.15e-05
.param mcm5m2_cc_w_4_000_s_10_000=1.21e-11
.param mcm5m2_cf_w_4_000_s_10_000=3.29e-11
.param mcm5m2_ca_w_4_000_s_12_000=1.15e-05
.param mcm5m2_cc_w_4_000_s_12_000=9.55e-12
.param mcm5m2_cf_w_4_000_s_12_000=3.52e-11
.param mcm5m3_ca_w_1_600_s_1_600=1.99e-05
.param mcm5m3_cc_w_1_600_s_1_600=6.33e-11
.param mcm5m3_cf_w_1_600_s_1_600=1.42e-11
.param mcm5m3_ca_w_1_600_s_1_700=1.99e-05
.param mcm5m3_cc_w_1_600_s_1_700=5.96e-11
.param mcm5m3_cf_w_1_600_s_1_700=1.50e-11
.param mcm5m3_ca_w_1_600_s_1_900=1.99e-05
.param mcm5m3_cc_w_1_600_s_1_900=5.33e-11
.param mcm5m3_cf_w_1_600_s_1_900=1.65e-11
.param mcm5m3_ca_w_1_600_s_2_000=1.99e-05
.param mcm5m3_cc_w_1_600_s_2_000=5.06e-11
.param mcm5m3_cf_w_1_600_s_2_000=1.72e-11
.param mcm5m3_ca_w_1_600_s_2_400=1.99e-05
.param mcm5m3_cc_w_1_600_s_2_400=4.21e-11
.param mcm5m3_cf_w_1_600_s_2_400=2.00e-11
.param mcm5m3_ca_w_1_600_s_2_800=1.99e-05
.param mcm5m3_cc_w_1_600_s_2_800=3.58e-11
.param mcm5m3_cf_w_1_600_s_2_800=2.25e-11
.param mcm5m3_ca_w_1_600_s_3_200=1.99e-05
.param mcm5m3_cc_w_1_600_s_3_200=3.11e-11
.param mcm5m3_cf_w_1_600_s_3_200=2.48e-11
.param mcm5m3_ca_w_1_600_s_4_800=1.99e-05
.param mcm5m3_cc_w_1_600_s_4_800=1.94e-11
.param mcm5m3_cf_w_1_600_s_4_800=3.19e-11
.param mcm5m3_ca_w_1_600_s_10_000=1.99e-05
.param mcm5m3_cc_w_1_600_s_10_000=6.90e-12
.param mcm5m3_cf_w_1_600_s_10_000=4.24e-11
.param mcm5m3_ca_w_1_600_s_12_000=1.99e-05
.param mcm5m3_cc_w_1_600_s_12_000=5.20e-12
.param mcm5m3_cf_w_1_600_s_12_000=4.41e-11
.param mcm5m3_ca_w_4_000_s_1_600=1.99e-05
.param mcm5m3_cc_w_4_000_s_1_600=6.86e-11
.param mcm5m3_cf_w_4_000_s_1_600=1.42e-11
.param mcm5m3_ca_w_4_000_s_1_700=1.99e-05
.param mcm5m3_cc_w_4_000_s_1_700=6.48e-11
.param mcm5m3_cf_w_4_000_s_1_700=1.50e-11
.param mcm5m3_ca_w_4_000_s_1_900=1.99e-05
.param mcm5m3_cc_w_4_000_s_1_900=5.83e-11
.param mcm5m3_cf_w_4_000_s_1_900=1.65e-11
.param mcm5m3_ca_w_4_000_s_2_000=1.99e-05
.param mcm5m3_cc_w_4_000_s_2_000=5.55e-11
.param mcm5m3_cf_w_4_000_s_2_000=1.72e-11
.param mcm5m3_ca_w_4_000_s_2_400=1.99e-05
.param mcm5m3_cc_w_4_000_s_2_400=4.66e-11
.param mcm5m3_cf_w_4_000_s_2_400=2.00e-11
.param mcm5m3_ca_w_4_000_s_2_800=1.99e-05
.param mcm5m3_cc_w_4_000_s_2_800=4.01e-11
.param mcm5m3_cf_w_4_000_s_2_800=2.25e-11
.param mcm5m3_ca_w_4_000_s_3_200=1.99e-05
.param mcm5m3_cc_w_4_000_s_3_200=3.52e-11
.param mcm5m3_cf_w_4_000_s_3_200=2.48e-11
.param mcm5m3_ca_w_4_000_s_4_800=1.99e-05
.param mcm5m3_cc_w_4_000_s_4_800=2.30e-11
.param mcm5m3_cf_w_4_000_s_4_800=3.21e-11
.param mcm5m3_ca_w_4_000_s_10_000=1.99e-05
.param mcm5m3_cc_w_4_000_s_10_000=9.15e-12
.param mcm5m3_cf_w_4_000_s_10_000=4.33e-11
.param mcm5m3_ca_w_4_000_s_12_000=1.99e-05
.param mcm5m3_cc_w_4_000_s_12_000=7.10e-12
.param mcm5m3_cf_w_4_000_s_12_000=4.53e-11
.param mcm5m4_ca_w_1_600_s_1_600=6.84e-05
.param mcm5m4_cc_w_1_600_s_1_600=5.05e-11
.param mcm5m4_cf_w_1_600_s_1_600=3.82e-11
.param mcm5m4_ca_w_1_600_s_1_700=6.84e-05
.param mcm5m4_cc_w_1_600_s_1_700=4.69e-11
.param mcm5m4_cf_w_1_600_s_1_700=3.97e-11
.param mcm5m4_ca_w_1_600_s_1_900=6.84e-05
.param mcm5m4_cc_w_1_600_s_1_900=4.09e-11
.param mcm5m4_cf_w_1_600_s_1_900=4.24e-11
.param mcm5m4_ca_w_1_600_s_2_000=6.84e-05
.param mcm5m4_cc_w_1_600_s_2_000=3.84e-11
.param mcm5m4_cf_w_1_600_s_2_000=4.37e-11
.param mcm5m4_ca_w_1_600_s_2_400=6.84e-05
.param mcm5m4_cc_w_1_600_s_2_400=3.06e-11
.param mcm5m4_cf_w_1_600_s_2_400=4.81e-11
.param mcm5m4_ca_w_1_600_s_2_800=6.84e-05
.param mcm5m4_cc_w_1_600_s_2_800=2.51e-11
.param mcm5m4_cf_w_1_600_s_2_800=5.17e-11
.param mcm5m4_ca_w_1_600_s_3_200=6.84e-05
.param mcm5m4_cc_w_1_600_s_3_200=2.11e-11
.param mcm5m4_cf_w_1_600_s_3_200=5.45e-11
.param mcm5m4_ca_w_1_600_s_4_800=6.84e-05
.param mcm5m4_cc_w_1_600_s_4_800=1.20e-11
.param mcm5m4_cf_w_1_600_s_4_800=6.19e-11
.param mcm5m4_ca_w_1_600_s_10_000=6.84e-05
.param mcm5m4_cc_w_1_600_s_10_000=4.00e-12
.param mcm5m4_cf_w_1_600_s_10_000=6.96e-11
.param mcm5m4_ca_w_1_600_s_12_000=6.84e-05
.param mcm5m4_cc_w_1_600_s_12_000=2.95e-12
.param mcm5m4_cf_w_1_600_s_12_000=7.06e-11
.param mcm5m4_ca_w_4_000_s_1_600=6.84e-05
.param mcm5m4_cc_w_4_000_s_1_600=5.57e-11
.param mcm5m4_cf_w_4_000_s_1_600=3.82e-11
.param mcm5m4_ca_w_4_000_s_1_700=6.84e-05
.param mcm5m4_cc_w_4_000_s_1_700=5.21e-11
.param mcm5m4_cf_w_4_000_s_1_700=3.97e-11
.param mcm5m4_ca_w_4_000_s_1_900=6.84e-05
.param mcm5m4_cc_w_4_000_s_1_900=4.59e-11
.param mcm5m4_cf_w_4_000_s_1_900=4.24e-11
.param mcm5m4_ca_w_4_000_s_2_000=6.84e-05
.param mcm5m4_cc_w_4_000_s_2_000=4.33e-11
.param mcm5m4_cf_w_4_000_s_2_000=4.37e-11
.param mcm5m4_ca_w_4_000_s_2_400=6.84e-05
.param mcm5m4_cc_w_4_000_s_2_400=3.52e-11
.param mcm5m4_cf_w_4_000_s_2_400=4.82e-11
.param mcm5m4_ca_w_4_000_s_2_800=6.84e-05
.param mcm5m4_cc_w_4_000_s_2_800=2.95e-11
.param mcm5m4_cf_w_4_000_s_2_800=5.17e-11
.param mcm5m4_ca_w_4_000_s_3_200=6.84e-05
.param mcm5m4_cc_w_4_000_s_3_200=2.52e-11
.param mcm5m4_cf_w_4_000_s_3_200=5.46e-11
.param mcm5m4_ca_w_4_000_s_4_800=6.84e-05
.param mcm5m4_cc_w_4_000_s_4_800=1.56e-11
.param mcm5m4_cf_w_4_000_s_4_800=6.23e-11
.param mcm5m4_ca_w_4_000_s_10_000=6.84e-05
.param mcm5m4_cc_w_4_000_s_10_000=6.00e-12
.param mcm5m4_cf_w_4_000_s_10_000=7.12e-11
.param mcm5m4_ca_w_4_000_s_12_000=6.84e-05
.param mcm5m4_cc_w_4_000_s_12_000=4.60e-12
.param mcm5m4_cf_w_4_000_s_12_000=7.26e-11
.param mcrdlf_ca_w_10_000_s_5_000=2.57e-06
.param mcrdlf_cc_w_10_000_s_5_000=5.16e-11
.param mcrdlf_cf_w_10_000_s_5_000=5.97e-12
.param mcrdlf_ca_w_10_000_s_8_000=2.57e-06
.param mcrdlf_cc_w_10_000_s_8_000=3.75e-11
.param mcrdlf_cf_w_10_000_s_8_000=9.04e-12
.param mcrdlf_ca_w_10_000_s_10_000=2.57e-06
.param mcrdlf_cc_w_10_000_s_10_000=3.20e-11
.param mcrdlf_cf_w_10_000_s_10_000=1.09e-11
.param mcrdlf_ca_w_10_000_s_12_000=2.57e-06
.param mcrdlf_cc_w_10_000_s_12_000=2.80e-11
.param mcrdlf_cf_w_10_000_s_12_000=1.26e-11
.param mcrdlf_ca_w_10_000_s_30_000=2.57e-06
.param mcrdlf_cc_w_10_000_s_30_000=1.23e-11
.param mcrdlf_cf_w_10_000_s_30_000=2.28e-11
.param mcrdlf_ca_w_40_000_s_5_000=2.57e-06
.param mcrdlf_cc_w_40_000_s_5_000=6.29e-11
.param mcrdlf_cf_w_40_000_s_5_000=6.08e-12
.param mcrdlf_ca_w_40_000_s_8_000=2.57e-06
.param mcrdlf_cc_w_40_000_s_8_000=4.79e-11
.param mcrdlf_cf_w_40_000_s_8_000=9.16e-12
.param mcrdlf_ca_w_40_000_s_10_000=2.57e-06
.param mcrdlf_cc_w_40_000_s_10_000=4.20e-11
.param mcrdlf_cf_w_40_000_s_10_000=1.10e-11
.param mcrdlf_ca_w_40_000_s_12_000=2.57e-06
.param mcrdlf_cc_w_40_000_s_12_000=3.74e-11
.param mcrdlf_cf_w_40_000_s_12_000=1.27e-11
.param mcrdlf_ca_w_40_000_s_30_000=2.57e-06
.param mcrdlf_cc_w_40_000_s_30_000=1.95e-11
.param mcrdlf_cf_w_40_000_s_30_000=2.35e-11
.param mcrdld_ca_w_10_000_s_5_000=2.63e-06
.param mcrdld_cc_w_10_000_s_5_000=5.14e-11
.param mcrdld_cf_w_10_000_s_5_000=6.11e-12
.param mcrdld_ca_w_10_000_s_8_000=2.63e-06
.param mcrdld_cc_w_10_000_s_8_000=3.73e-11
.param mcrdld_cf_w_10_000_s_8_000=9.23e-12
.param mcrdld_ca_w_10_000_s_10_000=2.63e-06
.param mcrdld_cc_w_10_000_s_10_000=3.18e-11
.param mcrdld_cf_w_10_000_s_10_000=1.11e-11
.param mcrdld_ca_w_10_000_s_12_000=2.63e-06
.param mcrdld_cc_w_10_000_s_12_000=2.78e-11
.param mcrdld_cf_w_10_000_s_12_000=1.28e-11
.param mcrdld_ca_w_10_000_s_30_000=2.63e-06
.param mcrdld_cc_w_10_000_s_30_000=1.22e-11
.param mcrdld_cf_w_10_000_s_30_000=2.31e-11
.param mcrdld_ca_w_40_000_s_5_000=2.63e-06
.param mcrdld_cc_w_40_000_s_5_000=6.27e-11
.param mcrdld_cf_w_40_000_s_5_000=6.23e-12
.param mcrdld_ca_w_40_000_s_8_000=2.63e-06
.param mcrdld_cc_w_40_000_s_8_000=4.76e-11
.param mcrdld_cf_w_40_000_s_8_000=9.36e-12
.param mcrdld_ca_w_40_000_s_10_000=2.63e-06
.param mcrdld_cc_w_40_000_s_10_000=4.17e-11
.param mcrdld_cf_w_40_000_s_10_000=1.12e-11
.param mcrdld_ca_w_40_000_s_12_000=2.63e-06
.param mcrdld_cc_w_40_000_s_12_000=3.72e-11
.param mcrdld_cf_w_40_000_s_12_000=1.30e-11
.param mcrdld_ca_w_40_000_s_30_000=2.63e-06
.param mcrdld_cc_w_40_000_s_30_000=1.94e-11
.param mcrdld_cf_w_40_000_s_30_000=2.38e-11
.param mcrdlp1_ca_w_10_000_s_5_000=2.68e-06
.param mcrdlp1_cc_w_10_000_s_5_000=5.12e-11
.param mcrdlp1_cf_w_10_000_s_5_000=6.21e-12
.param mcrdlp1_ca_w_10_000_s_8_000=2.68e-06
.param mcrdlp1_cc_w_10_000_s_8_000=3.71e-11
.param mcrdlp1_cf_w_10_000_s_8_000=9.38e-12
.param mcrdlp1_ca_w_10_000_s_10_000=2.68e-06
.param mcrdlp1_cc_w_10_000_s_10_000=3.16e-11
.param mcrdlp1_cf_w_10_000_s_10_000=1.13e-11
.param mcrdlp1_ca_w_10_000_s_12_000=2.68e-06
.param mcrdlp1_cc_w_10_000_s_12_000=2.76e-11
.param mcrdlp1_cf_w_10_000_s_12_000=1.31e-11
.param mcrdlp1_ca_w_10_000_s_30_000=2.68e-06
.param mcrdlp1_cc_w_10_000_s_30_000=1.21e-11
.param mcrdlp1_cf_w_10_000_s_30_000=2.34e-11
.param mcrdlp1_ca_w_40_000_s_5_000=2.68e-06
.param mcrdlp1_cc_w_40_000_s_5_000=6.25e-11
.param mcrdlp1_cf_w_40_000_s_5_000=6.36e-12
.param mcrdlp1_ca_w_40_000_s_8_000=2.68e-06
.param mcrdlp1_cc_w_40_000_s_8_000=4.75e-11
.param mcrdlp1_cf_w_40_000_s_8_000=9.54e-12
.param mcrdlp1_ca_w_40_000_s_10_000=2.68e-06
.param mcrdlp1_cc_w_40_000_s_10_000=4.15e-11
.param mcrdlp1_cf_w_40_000_s_10_000=1.15e-11
.param mcrdlp1_ca_w_40_000_s_12_000=2.68e-06
.param mcrdlp1_cc_w_40_000_s_12_000=3.71e-11
.param mcrdlp1_cf_w_40_000_s_12_000=1.32e-11
.param mcrdlp1_ca_w_40_000_s_30_000=2.68e-06
.param mcrdlp1_cc_w_40_000_s_30_000=1.92e-11
.param mcrdlp1_cf_w_40_000_s_30_000=2.41e-11
.param mcrdll1_ca_w_10_000_s_5_000=2.78e-06
.param mcrdll1_cc_w_10_000_s_5_000=5.09e-11
.param mcrdll1_cf_w_10_000_s_5_000=6.41e-12
.param mcrdll1_ca_w_10_000_s_8_000=2.78e-06
.param mcrdll1_cc_w_10_000_s_8_000=3.68e-11
.param mcrdll1_cf_w_10_000_s_8_000=9.67e-12
.param mcrdll1_ca_w_10_000_s_10_000=2.78e-06
.param mcrdll1_cc_w_10_000_s_10_000=3.13e-11
.param mcrdll1_cf_w_10_000_s_10_000=1.16e-11
.param mcrdll1_ca_w_10_000_s_12_000=2.78e-06
.param mcrdll1_cc_w_10_000_s_12_000=2.74e-11
.param mcrdll1_cf_w_10_000_s_12_000=1.34e-11
.param mcrdll1_ca_w_10_000_s_30_000=2.78e-06
.param mcrdll1_cc_w_10_000_s_30_000=1.18e-11
.param mcrdll1_cf_w_10_000_s_30_000=2.38e-11
.param mcrdll1_ca_w_40_000_s_5_000=2.78e-06
.param mcrdll1_cc_w_40_000_s_5_000=6.22e-11
.param mcrdll1_cf_w_40_000_s_5_000=6.49e-12
.param mcrdll1_ca_w_40_000_s_8_000=2.78e-06
.param mcrdll1_cc_w_40_000_s_8_000=4.72e-11
.param mcrdll1_cf_w_40_000_s_8_000=9.76e-12
.param mcrdll1_ca_w_40_000_s_10_000=2.78e-06
.param mcrdll1_cc_w_40_000_s_10_000=4.12e-11
.param mcrdll1_cf_w_40_000_s_10_000=1.17e-11
.param mcrdll1_ca_w_40_000_s_12_000=2.78e-06
.param mcrdll1_cc_w_40_000_s_12_000=3.68e-11
.param mcrdll1_cf_w_40_000_s_12_000=1.35e-11
.param mcrdll1_ca_w_40_000_s_30_000=2.78e-06
.param mcrdll1_cc_w_40_000_s_30_000=1.90e-11
.param mcrdll1_cf_w_40_000_s_30_000=2.45e-11
.param mcrdlm1_ca_w_10_000_s_5_000=2.93e-06
.param mcrdlm1_cc_w_10_000_s_5_000=5.04e-11
.param mcrdlm1_cf_w_10_000_s_5_000=6.73e-12
.param mcrdlm1_ca_w_10_000_s_8_000=2.93e-06
.param mcrdlm1_cc_w_10_000_s_8_000=3.63e-11
.param mcrdlm1_cf_w_10_000_s_8_000=1.01e-11
.param mcrdlm1_ca_w_10_000_s_10_000=2.93e-06
.param mcrdlm1_cc_w_10_000_s_10_000=3.09e-11
.param mcrdlm1_cf_w_10_000_s_10_000=1.21e-11
.param mcrdlm1_ca_w_10_000_s_12_000=2.93e-06
.param mcrdlm1_cc_w_10_000_s_12_000=2.69e-11
.param mcrdlm1_cf_w_10_000_s_12_000=1.40e-11
.param mcrdlm1_ca_w_10_000_s_30_000=2.93e-06
.param mcrdlm1_cc_w_10_000_s_30_000=1.15e-11
.param mcrdlm1_cf_w_10_000_s_30_000=2.45e-11
.param mcrdlm1_ca_w_40_000_s_5_000=2.93e-06
.param mcrdlm1_cc_w_40_000_s_5_000=6.17e-11
.param mcrdlm1_cf_w_40_000_s_5_000=6.82e-12
.param mcrdlm1_ca_w_40_000_s_8_000=2.93e-06
.param mcrdlm1_cc_w_40_000_s_8_000=4.67e-11
.param mcrdlm1_cf_w_40_000_s_8_000=1.02e-11
.param mcrdlm1_ca_w_40_000_s_10_000=2.93e-06
.param mcrdlm1_cc_w_40_000_s_10_000=4.08e-11
.param mcrdlm1_cf_w_40_000_s_10_000=1.22e-11
.param mcrdlm1_ca_w_40_000_s_12_000=2.93e-06
.param mcrdlm1_cc_w_40_000_s_12_000=3.64e-11
.param mcrdlm1_cf_w_40_000_s_12_000=1.41e-11
.param mcrdlm1_ca_w_40_000_s_30_000=2.93e-06
.param mcrdlm1_cc_w_40_000_s_30_000=1.86e-11
.param mcrdlm1_cf_w_40_000_s_30_000=2.53e-11
.param mcrdlm2_ca_w_10_000_s_5_000=3.10e-06
.param mcrdlm2_cc_w_10_000_s_5_000=4.99e-11
.param mcrdlm2_cf_w_10_000_s_5_000=7.07e-12
.param mcrdlm2_ca_w_10_000_s_8_000=3.10e-06
.param mcrdlm2_cc_w_10_000_s_8_000=3.59e-11
.param mcrdlm2_cf_w_10_000_s_8_000=1.06e-11
.param mcrdlm2_ca_w_10_000_s_10_000=3.10e-06
.param mcrdlm2_cc_w_10_000_s_10_000=3.04e-11
.param mcrdlm2_cf_w_10_000_s_10_000=1.27e-11
.param mcrdlm2_ca_w_10_000_s_12_000=3.10e-06
.param mcrdlm2_cc_w_10_000_s_12_000=2.65e-11
.param mcrdlm2_cf_w_10_000_s_12_000=1.46e-11
.param mcrdlm2_ca_w_10_000_s_30_000=3.10e-06
.param mcrdlm2_cc_w_10_000_s_30_000=1.12e-11
.param mcrdlm2_cf_w_10_000_s_30_000=2.52e-11
.param mcrdlm2_ca_w_40_000_s_5_000=3.10e-06
.param mcrdlm2_cc_w_40_000_s_5_000=6.12e-11
.param mcrdlm2_cf_w_40_000_s_5_000=7.14e-12
.param mcrdlm2_ca_w_40_000_s_8_000=3.10e-06
.param mcrdlm2_cc_w_40_000_s_8_000=4.62e-11
.param mcrdlm2_cf_w_40_000_s_8_000=1.07e-11
.param mcrdlm2_ca_w_40_000_s_10_000=3.10e-06
.param mcrdlm2_cc_w_40_000_s_10_000=4.03e-11
.param mcrdlm2_cf_w_40_000_s_10_000=1.28e-11
.param mcrdlm2_ca_w_40_000_s_12_000=3.10e-06
.param mcrdlm2_cc_w_40_000_s_12_000=3.58e-11
.param mcrdlm2_cf_w_40_000_s_12_000=1.47e-11
.param mcrdlm2_ca_w_40_000_s_30_000=3.10e-06
.param mcrdlm2_cc_w_40_000_s_30_000=1.83e-11
.param mcrdlm2_cf_w_40_000_s_30_000=2.60e-11
.param mcrdlm3_ca_w_10_000_s_5_000=3.50e-06
.param mcrdlm3_cc_w_10_000_s_5_000=4.89e-11
.param mcrdlm3_cf_w_10_000_s_5_000=7.87e-12
.param mcrdlm3_ca_w_10_000_s_8_000=3.50e-06
.param mcrdlm3_cc_w_10_000_s_8_000=3.49e-11
.param mcrdlm3_cf_w_10_000_s_8_000=1.17e-11
.param mcrdlm3_ca_w_10_000_s_10_000=3.50e-06
.param mcrdlm3_cc_w_10_000_s_10_000=2.95e-11
.param mcrdlm3_cf_w_10_000_s_10_000=1.39e-11
.param mcrdlm3_ca_w_10_000_s_12_000=3.50e-06
.param mcrdlm3_cc_w_10_000_s_12_000=2.55e-11
.param mcrdlm3_cf_w_10_000_s_12_000=1.59e-11
.param mcrdlm3_ca_w_10_000_s_30_000=3.50e-06
.param mcrdlm3_cc_w_10_000_s_30_000=1.06e-11
.param mcrdlm3_cf_w_10_000_s_30_000=2.67e-11
.param mcrdlm3_ca_w_40_000_s_5_000=3.50e-06
.param mcrdlm3_cc_w_40_000_s_5_000=6.02e-11
.param mcrdlm3_cf_w_40_000_s_5_000=7.93e-12
.param mcrdlm3_ca_w_40_000_s_8_000=3.50e-06
.param mcrdlm3_cc_w_40_000_s_8_000=4.52e-11
.param mcrdlm3_cf_w_40_000_s_8_000=1.18e-11
.param mcrdlm3_ca_w_40_000_s_10_000=3.50e-06
.param mcrdlm3_cc_w_40_000_s_10_000=3.93e-11
.param mcrdlm3_cf_w_40_000_s_10_000=1.40e-11
.param mcrdlm3_ca_w_40_000_s_12_000=3.50e-06
.param mcrdlm3_cc_w_40_000_s_12_000=3.50e-11
.param mcrdlm3_cf_w_40_000_s_12_000=1.60e-11
.param mcrdlm3_ca_w_40_000_s_30_000=3.50e-06
.param mcrdlm3_cc_w_40_000_s_30_000=1.77e-11
.param mcrdlm3_cf_w_40_000_s_30_000=2.77e-11
.param mcrdlm4_ca_w_10_000_s_5_000=4.00e-06
.param mcrdlm4_cc_w_10_000_s_5_000=4.78e-11
.param mcrdlm4_cf_w_10_000_s_5_000=8.79e-12
.param mcrdlm4_ca_w_10_000_s_8_000=4.00e-06
.param mcrdlm4_cc_w_10_000_s_8_000=3.38e-11
.param mcrdlm4_cf_w_10_000_s_8_000=1.30e-11
.param mcrdlm4_ca_w_10_000_s_10_000=4.00e-06
.param mcrdlm4_cc_w_10_000_s_10_000=2.85e-11
.param mcrdlm4_cf_w_10_000_s_10_000=1.54e-11
.param mcrdlm4_ca_w_10_000_s_12_000=4.00e-06
.param mcrdlm4_cc_w_10_000_s_12_000=2.45e-11
.param mcrdlm4_cf_w_10_000_s_12_000=1.75e-11
.param mcrdlm4_ca_w_10_000_s_30_000=4.00e-06
.param mcrdlm4_cc_w_10_000_s_30_000=9.97e-12
.param mcrdlm4_cf_w_10_000_s_30_000=2.84e-11
.param mcrdlm4_ca_w_40_000_s_5_000=4.00e-06
.param mcrdlm4_cc_w_40_000_s_5_000=5.90e-11
.param mcrdlm4_cf_w_40_000_s_5_000=8.71e-12
.param mcrdlm4_ca_w_40_000_s_8_000=4.00e-06
.param mcrdlm4_cc_w_40_000_s_8_000=4.41e-11
.param mcrdlm4_cf_w_40_000_s_8_000=1.29e-11
.param mcrdlm4_ca_w_40_000_s_10_000=4.00e-06
.param mcrdlm4_cc_w_40_000_s_10_000=3.83e-11
.param mcrdlm4_cf_w_40_000_s_10_000=1.53e-11
.param mcrdlm4_ca_w_40_000_s_12_000=4.00e-06
.param mcrdlm4_cc_w_40_000_s_12_000=3.40e-11
.param mcrdlm4_cf_w_40_000_s_12_000=1.75e-11
.param mcrdlm4_ca_w_40_000_s_30_000=4.00e-06
.param mcrdlm4_cc_w_40_000_s_30_000=1.70e-11
.param mcrdlm4_cf_w_40_000_s_30_000=2.94e-11
.param mcrdlm5_ca_w_10_000_s_5_000=5.44e-06
.param mcrdlm5_cc_w_10_000_s_5_000=4.54e-11
.param mcrdlm5_cf_w_10_000_s_5_000=1.14e-11
.param mcrdlm5_ca_w_10_000_s_8_000=5.44e-06
.param mcrdlm5_cc_w_10_000_s_8_000=3.16e-11
.param mcrdlm5_cf_w_10_000_s_8_000=1.64e-11
.param mcrdlm5_ca_w_10_000_s_10_000=5.44e-06
.param mcrdlm5_cc_w_10_000_s_10_000=2.63e-11
.param mcrdlm5_cf_w_10_000_s_10_000=1.92e-11
.param mcrdlm5_ca_w_10_000_s_12_000=5.44e-06
.param mcrdlm5_cc_w_10_000_s_12_000=2.25e-11
.param mcrdlm5_cf_w_10_000_s_12_000=2.15e-11
.param mcrdlm5_ca_w_10_000_s_30_000=5.44e-06
.param mcrdlm5_cc_w_10_000_s_30_000=8.70e-12
.param mcrdlm5_cf_w_10_000_s_30_000=3.26e-11
.param mcrdlm5_ca_w_40_000_s_5_000=5.44e-06
.param mcrdlm5_cc_w_40_000_s_5_000=5.67e-11
.param mcrdlm5_cf_w_40_000_s_5_000=1.14e-11
.param mcrdlm5_ca_w_40_000_s_8_000=5.44e-06
.param mcrdlm5_cc_w_40_000_s_8_000=4.19e-11
.param mcrdlm5_cf_w_40_000_s_8_000=1.64e-11
.param mcrdlm5_ca_w_40_000_s_10_000=5.44e-06
.param mcrdlm5_cc_w_40_000_s_10_000=3.62e-11
.param mcrdlm5_cf_w_40_000_s_10_000=1.92e-11
.param mcrdlm5_ca_w_40_000_s_12_000=5.44e-06
.param mcrdlm5_cc_w_40_000_s_12_000=3.20e-11
.param mcrdlm5_cf_w_40_000_s_12_000=2.16e-11
.param mcrdlm5_ca_w_40_000_s_30_000=5.44e-06
.param mcrdlm5_cc_w_40_000_s_30_000=1.57e-11
.param mcrdlm5_cf_w_40_000_s_30_000=3.38e-11
.param mcl1p1f_ca_w_0_150_s_0_210=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_210=6.42e-11
.param mcl1p1f_cf_w_0_150_s_0_210=1.91e-11
.param mcl1p1f_ca_w_0_150_s_0_263=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_263=4.90e-11
.param mcl1p1f_cf_w_0_150_s_0_263=2.32e-11
.param mcl1p1f_ca_w_0_150_s_0_315=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_315=3.87e-11
.param mcl1p1f_cf_w_0_150_s_0_315=2.68e-11
.param mcl1p1f_ca_w_0_150_s_0_420=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_420=2.56e-11
.param mcl1p1f_cf_w_0_150_s_0_420=3.33e-11
.param mcl1p1f_ca_w_0_150_s_0_525=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_525=1.74e-11
.param mcl1p1f_cf_w_0_150_s_0_525=3.84e-11
.param mcl1p1f_ca_w_0_150_s_0_630=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_630=1.21e-11
.param mcl1p1f_cf_w_0_150_s_0_630=4.23e-11
.param mcl1p1f_ca_w_0_150_s_0_840=2.00e-04
.param mcl1p1f_cc_w_0_150_s_0_840=5.89e-12
.param mcl1p1f_cf_w_0_150_s_0_840=4.74e-11
.param mcl1p1f_ca_w_0_150_s_1_260=2.00e-04
.param mcl1p1f_cc_w_0_150_s_1_260=1.52e-12
.param mcl1p1f_cf_w_0_150_s_1_260=5.15e-11
.param mcl1p1f_ca_w_0_150_s_2_310=2.00e-04
.param mcl1p1f_cc_w_0_150_s_2_310=1.10e-13
.param mcl1p1f_cf_w_0_150_s_2_310=5.29e-11
.param mcl1p1f_ca_w_0_150_s_5_250=2.00e-04
.param mcl1p1f_cc_w_0_150_s_5_250=5.00e-15
.param mcl1p1f_cf_w_0_150_s_5_250=5.30e-11
.param mcl1p1f_ca_w_1_200_s_0_210=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_210=6.64e-11
.param mcl1p1f_cf_w_1_200_s_0_210=1.90e-11
.param mcl1p1f_ca_w_1_200_s_0_263=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_263=5.07e-11
.param mcl1p1f_cf_w_1_200_s_0_263=2.31e-11
.param mcl1p1f_ca_w_1_200_s_0_315=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_315=4.02e-11
.param mcl1p1f_cf_w_1_200_s_0_315=2.69e-11
.param mcl1p1f_ca_w_1_200_s_0_420=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_420=2.66e-11
.param mcl1p1f_cf_w_1_200_s_0_420=3.34e-11
.param mcl1p1f_ca_w_1_200_s_0_525=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_525=1.81e-11
.param mcl1p1f_cf_w_1_200_s_0_525=3.86e-11
.param mcl1p1f_ca_w_1_200_s_0_630=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_630=1.26e-11
.param mcl1p1f_cf_w_1_200_s_0_630=4.26e-11
.param mcl1p1f_ca_w_1_200_s_0_840=2.00e-04
.param mcl1p1f_cc_w_1_200_s_0_840=6.20e-12
.param mcl1p1f_cf_w_1_200_s_0_840=4.80e-11
.param mcl1p1f_ca_w_1_200_s_1_260=2.00e-04
.param mcl1p1f_cc_w_1_200_s_1_260=1.60e-12
.param mcl1p1f_cf_w_1_200_s_1_260=5.23e-11
.param mcl1p1f_ca_w_1_200_s_2_310=2.00e-04
.param mcl1p1f_cc_w_1_200_s_2_310=1.50e-13
.param mcl1p1f_cf_w_1_200_s_2_310=5.37e-11
.param mcl1p1f_ca_w_1_200_s_5_250=2.00e-04
.param mcl1p1f_cc_w_1_200_s_5_250=0.00e+00
.param mcl1p1f_cf_w_1_200_s_5_250=5.38e-11
.param mcm1p1f_ca_w_0_150_s_0_210=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_210=6.98e-11
.param mcm1p1f_cf_w_0_150_s_0_210=1.48e-11
.param mcm1p1f_ca_w_0_150_s_0_263=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_263=5.50e-11
.param mcm1p1f_cf_w_0_150_s_0_263=1.80e-11
.param mcm1p1f_ca_w_0_150_s_0_315=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_315=4.48e-11
.param mcm1p1f_cf_w_0_150_s_0_315=2.09e-11
.param mcm1p1f_ca_w_0_150_s_0_420=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_420=3.17e-11
.param mcm1p1f_cf_w_0_150_s_0_420=2.64e-11
.param mcm1p1f_ca_w_0_150_s_0_525=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_525=2.33e-11
.param mcm1p1f_cf_w_0_150_s_0_525=3.09e-11
.param mcm1p1f_ca_w_0_150_s_0_630=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_630=1.75e-11
.param mcm1p1f_cf_w_0_150_s_0_630=3.45e-11
.param mcm1p1f_ca_w_0_150_s_0_840=1.51e-04
.param mcm1p1f_cc_w_0_150_s_0_840=1.03e-11
.param mcm1p1f_cf_w_0_150_s_0_840=4.00e-11
.param mcm1p1f_ca_w_0_150_s_1_260=1.51e-04
.param mcm1p1f_cc_w_0_150_s_1_260=3.78e-12
.param mcm1p1f_cf_w_0_150_s_1_260=4.57e-11
.param mcm1p1f_ca_w_0_150_s_2_310=1.51e-04
.param mcm1p1f_cc_w_0_150_s_2_310=3.70e-13
.param mcm1p1f_cf_w_0_150_s_2_310=4.88e-11
.param mcm1p1f_ca_w_0_150_s_5_250=1.51e-04
.param mcm1p1f_cc_w_0_150_s_5_250=4.00e-14
.param mcm1p1f_cf_w_0_150_s_5_250=4.92e-11
.param mcm1p1f_ca_w_1_200_s_0_210=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_210=7.52e-11
.param mcm1p1f_cf_w_1_200_s_0_210=1.47e-11
.param mcm1p1f_ca_w_1_200_s_0_263=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_263=5.93e-11
.param mcm1p1f_cf_w_1_200_s_0_263=1.79e-11
.param mcm1p1f_ca_w_1_200_s_0_315=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_315=4.87e-11
.param mcm1p1f_cf_w_1_200_s_0_315=2.09e-11
.param mcm1p1f_ca_w_1_200_s_0_420=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_420=3.46e-11
.param mcm1p1f_cf_w_1_200_s_0_420=2.64e-11
.param mcm1p1f_ca_w_1_200_s_0_525=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_525=2.57e-11
.param mcm1p1f_cf_w_1_200_s_0_525=3.11e-11
.param mcm1p1f_ca_w_1_200_s_0_630=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_630=1.95e-11
.param mcm1p1f_cf_w_1_200_s_0_630=3.49e-11
.param mcm1p1f_ca_w_1_200_s_0_840=1.51e-04
.param mcm1p1f_cc_w_1_200_s_0_840=1.16e-11
.param mcm1p1f_cf_w_1_200_s_0_840=4.07e-11
.param mcm1p1f_ca_w_1_200_s_1_260=1.51e-04
.param mcm1p1f_cc_w_1_200_s_1_260=4.37e-12
.param mcm1p1f_cf_w_1_200_s_1_260=4.70e-11
.param mcm1p1f_ca_w_1_200_s_2_310=1.51e-04
.param mcm1p1f_cc_w_1_200_s_2_310=4.60e-13
.param mcm1p1f_cf_w_1_200_s_2_310=5.07e-11
.param mcm1p1f_ca_w_1_200_s_5_250=1.51e-04
.param mcm1p1f_cc_w_1_200_s_5_250=0.00e+00
.param mcm1p1f_cf_w_1_200_s_5_250=5.11e-11
.param mcm2p1f_ca_w_0_150_s_0_210=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_210=7.25e-11
.param mcm2p1f_cf_w_0_150_s_0_210=1.28e-11
.param mcm2p1f_ca_w_0_150_s_0_263=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_263=5.80e-11
.param mcm2p1f_cf_w_0_150_s_0_263=1.56e-11
.param mcm2p1f_ca_w_0_150_s_0_315=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_315=4.81e-11
.param mcm2p1f_cf_w_0_150_s_0_315=1.82e-11
.param mcm2p1f_ca_w_0_150_s_0_420=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_420=3.53e-11
.param mcm2p1f_cf_w_0_150_s_0_420=2.30e-11
.param mcm2p1f_ca_w_0_150_s_0_525=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_525=2.71e-11
.param mcm2p1f_cf_w_0_150_s_0_525=2.71e-11
.param mcm2p1f_ca_w_0_150_s_0_630=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_630=2.13e-11
.param mcm2p1f_cf_w_0_150_s_0_630=3.05e-11
.param mcm2p1f_ca_w_0_150_s_0_840=1.31e-04
.param mcm2p1f_cc_w_0_150_s_0_840=1.37e-11
.param mcm2p1f_cf_w_0_150_s_0_840=3.58e-11
.param mcm2p1f_ca_w_0_150_s_1_260=1.31e-04
.param mcm2p1f_cc_w_0_150_s_1_260=6.29e-12
.param mcm2p1f_cf_w_0_150_s_1_260=4.20e-11
.param mcm2p1f_ca_w_0_150_s_2_310=1.31e-04
.param mcm2p1f_cc_w_0_150_s_2_310=1.12e-12
.param mcm2p1f_cf_w_0_150_s_2_310=4.67e-11
.param mcm2p1f_ca_w_0_150_s_5_250=1.31e-04
.param mcm2p1f_cc_w_0_150_s_5_250=5.00e-14
.param mcm2p1f_cf_w_0_150_s_5_250=4.78e-11
.param mcm2p1f_ca_w_1_200_s_0_210=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_210=8.17e-11
.param mcm2p1f_cf_w_1_200_s_0_210=1.27e-11
.param mcm2p1f_ca_w_1_200_s_0_263=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_263=6.59e-11
.param mcm2p1f_cf_w_1_200_s_0_263=1.56e-11
.param mcm2p1f_ca_w_1_200_s_0_315=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_315=5.52e-11
.param mcm2p1f_cf_w_1_200_s_0_315=1.82e-11
.param mcm2p1f_ca_w_1_200_s_0_420=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_420=4.11e-11
.param mcm2p1f_cf_w_1_200_s_0_420=2.30e-11
.param mcm2p1f_ca_w_1_200_s_0_525=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_525=3.20e-11
.param mcm2p1f_cf_w_1_200_s_0_525=2.72e-11
.param mcm2p1f_ca_w_1_200_s_0_630=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_630=2.56e-11
.param mcm2p1f_cf_w_1_200_s_0_630=3.08e-11
.param mcm2p1f_ca_w_1_200_s_0_840=1.31e-04
.param mcm2p1f_cc_w_1_200_s_0_840=1.70e-11
.param mcm2p1f_cf_w_1_200_s_0_840=3.65e-11
.param mcm2p1f_ca_w_1_200_s_1_260=1.31e-04
.param mcm2p1f_cc_w_1_200_s_1_260=8.21e-12
.param mcm2p1f_cf_w_1_200_s_1_260=4.36e-11
.param mcm2p1f_ca_w_1_200_s_2_310=1.31e-04
.param mcm2p1f_cc_w_1_200_s_2_310=1.59e-12
.param mcm2p1f_cf_w_1_200_s_2_310=4.97e-11
.param mcm2p1f_ca_w_1_200_s_5_250=1.31e-04
.param mcm2p1f_cc_w_1_200_s_5_250=3.50e-14
.param mcm2p1f_cf_w_1_200_s_5_250=5.12e-11
.param mcm3p1f_ca_w_0_150_s_0_210=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_210=7.38e-11
.param mcm3p1f_cf_w_0_150_s_0_210=1.19e-11
.param mcm3p1f_ca_w_0_150_s_0_263=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_263=5.94e-11
.param mcm3p1f_cf_w_0_150_s_0_263=1.45e-11
.param mcm3p1f_ca_w_0_150_s_0_315=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_315=4.99e-11
.param mcm3p1f_cf_w_0_150_s_0_315=1.69e-11
.param mcm3p1f_ca_w_0_150_s_0_420=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_420=3.71e-11
.param mcm3p1f_cf_w_0_150_s_0_420=2.14e-11
.param mcm3p1f_ca_w_0_150_s_0_525=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_525=2.91e-11
.param mcm3p1f_cf_w_0_150_s_0_525=2.53e-11
.param mcm3p1f_ca_w_0_150_s_0_630=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_630=2.34e-11
.param mcm3p1f_cf_w_0_150_s_0_630=2.85e-11
.param mcm3p1f_ca_w_0_150_s_0_840=1.22e-04
.param mcm3p1f_cc_w_0_150_s_0_840=1.58e-11
.param mcm3p1f_cf_w_0_150_s_0_840=3.37e-11
.param mcm3p1f_ca_w_0_150_s_1_260=1.22e-04
.param mcm3p1f_cc_w_0_150_s_1_260=7.92e-12
.param mcm3p1f_cf_w_0_150_s_1_260=4.01e-11
.param mcm3p1f_ca_w_0_150_s_2_310=1.22e-04
.param mcm3p1f_cc_w_0_150_s_2_310=1.95e-12
.param mcm3p1f_cf_w_0_150_s_2_310=4.55e-11
.param mcm3p1f_ca_w_0_150_s_5_250=1.22e-04
.param mcm3p1f_cc_w_0_150_s_5_250=1.05e-13
.param mcm3p1f_cf_w_0_150_s_5_250=4.73e-11
.param mcm3p1f_ca_w_1_200_s_0_210=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_210=8.57e-11
.param mcm3p1f_cf_w_1_200_s_0_210=1.19e-11
.param mcm3p1f_ca_w_1_200_s_0_263=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_263=6.98e-11
.param mcm3p1f_cf_w_1_200_s_0_263=1.45e-11
.param mcm3p1f_ca_w_1_200_s_0_315=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_315=5.93e-11
.param mcm3p1f_cf_w_1_200_s_0_315=1.69e-11
.param mcm3p1f_ca_w_1_200_s_0_420=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_420=4.51e-11
.param mcm3p1f_cf_w_1_200_s_0_420=2.14e-11
.param mcm3p1f_ca_w_1_200_s_0_525=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_525=3.60e-11
.param mcm3p1f_cf_w_1_200_s_0_525=2.54e-11
.param mcm3p1f_ca_w_1_200_s_0_630=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_630=2.96e-11
.param mcm3p1f_cf_w_1_200_s_0_630=2.88e-11
.param mcm3p1f_ca_w_1_200_s_0_840=1.22e-04
.param mcm3p1f_cc_w_1_200_s_0_840=2.08e-11
.param mcm3p1f_cf_w_1_200_s_0_840=3.44e-11
.param mcm3p1f_ca_w_1_200_s_1_260=1.22e-04
.param mcm3p1f_cc_w_1_200_s_1_260=1.13e-11
.param mcm3p1f_cf_w_1_200_s_1_260=4.16e-11
.param mcm3p1f_ca_w_1_200_s_2_310=1.22e-04
.param mcm3p1f_cc_w_1_200_s_2_310=3.11e-12
.param mcm3p1f_cf_w_1_200_s_2_310=4.90e-11
.param mcm3p1f_ca_w_1_200_s_5_250=1.22e-04
.param mcm3p1f_cc_w_1_200_s_5_250=1.50e-13
.param mcm3p1f_cf_w_1_200_s_5_250=5.19e-11
.param mcm4p1f_ca_w_0_150_s_0_210=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_210=7.48e-11
.param mcm4p1f_cf_w_0_150_s_0_210=1.14e-11
.param mcm4p1f_ca_w_0_150_s_0_263=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_263=6.03e-11
.param mcm4p1f_cf_w_0_150_s_0_263=1.38e-11
.param mcm4p1f_ca_w_0_150_s_0_315=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_315=5.10e-11
.param mcm4p1f_cf_w_0_150_s_0_315=1.61e-11
.param mcm4p1f_ca_w_0_150_s_0_420=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_420=3.83e-11
.param mcm4p1f_cf_w_0_150_s_0_420=2.04e-11
.param mcm4p1f_ca_w_0_150_s_0_525=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_525=3.05e-11
.param mcm4p1f_cf_w_0_150_s_0_525=2.40e-11
.param mcm4p1f_ca_w_0_150_s_0_630=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_630=2.49e-11
.param mcm4p1f_cf_w_0_150_s_0_630=2.72e-11
.param mcm4p1f_ca_w_0_150_s_0_840=1.16e-04
.param mcm4p1f_cc_w_0_150_s_0_840=1.74e-11
.param mcm4p1f_cf_w_0_150_s_0_840=3.22e-11
.param mcm4p1f_ca_w_0_150_s_1_260=1.16e-04
.param mcm4p1f_cc_w_0_150_s_1_260=9.22e-12
.param mcm4p1f_cf_w_0_150_s_1_260=3.88e-11
.param mcm4p1f_ca_w_0_150_s_2_310=1.16e-04
.param mcm4p1f_cc_w_0_150_s_2_310=2.78e-12
.param mcm4p1f_cf_w_0_150_s_2_310=4.45e-11
.param mcm4p1f_ca_w_0_150_s_5_250=1.16e-04
.param mcm4p1f_cc_w_0_150_s_5_250=2.45e-13
.param mcm4p1f_cf_w_0_150_s_5_250=4.71e-11
.param mcm4p1f_ca_w_1_200_s_0_210=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_210=8.87e-11
.param mcm4p1f_cf_w_1_200_s_0_210=1.13e-11
.param mcm4p1f_ca_w_1_200_s_0_263=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_263=7.30e-11
.param mcm4p1f_cf_w_1_200_s_0_263=1.38e-11
.param mcm4p1f_ca_w_1_200_s_0_315=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_315=6.24e-11
.param mcm4p1f_cf_w_1_200_s_0_315=1.61e-11
.param mcm4p1f_ca_w_1_200_s_0_420=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_420=4.83e-11
.param mcm4p1f_cf_w_1_200_s_0_420=2.04e-11
.param mcm4p1f_ca_w_1_200_s_0_525=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_525=3.93e-11
.param mcm4p1f_cf_w_1_200_s_0_525=2.42e-11
.param mcm4p1f_ca_w_1_200_s_0_630=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_630=3.28e-11
.param mcm4p1f_cf_w_1_200_s_0_630=2.75e-11
.param mcm4p1f_ca_w_1_200_s_0_840=1.16e-04
.param mcm4p1f_cc_w_1_200_s_0_840=2.40e-11
.param mcm4p1f_cf_w_1_200_s_0_840=3.29e-11
.param mcm4p1f_ca_w_1_200_s_1_260=1.16e-04
.param mcm4p1f_cc_w_1_200_s_1_260=1.42e-11
.param mcm4p1f_cf_w_1_200_s_1_260=4.01e-11
.param mcm4p1f_ca_w_1_200_s_2_310=1.16e-04
.param mcm4p1f_cc_w_1_200_s_2_310=4.91e-12
.param mcm4p1f_cf_w_1_200_s_2_310=4.84e-11
.param mcm4p1f_ca_w_1_200_s_5_250=1.16e-04
.param mcm4p1f_cc_w_1_200_s_5_250=4.80e-13
.param mcm4p1f_cf_w_1_200_s_5_250=5.27e-11
.param mcm5p1f_ca_w_0_150_s_0_210=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_210=7.51e-11
.param mcm5p1f_cf_w_0_150_s_0_210=1.11e-11
.param mcm5p1f_ca_w_0_150_s_0_263=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_263=6.08e-11
.param mcm5p1f_cf_w_0_150_s_0_263=1.34e-11
.param mcm5p1f_ca_w_0_150_s_0_315=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_315=5.15e-11
.param mcm5p1f_cf_w_0_150_s_0_315=1.57e-11
.param mcm5p1f_ca_w_0_150_s_0_420=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_420=3.89e-11
.param mcm5p1f_cf_w_0_150_s_0_420=1.99e-11
.param mcm5p1f_ca_w_0_150_s_0_525=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_525=3.12e-11
.param mcm5p1f_cf_w_0_150_s_0_525=2.34e-11
.param mcm5p1f_ca_w_0_150_s_0_630=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_630=2.56e-11
.param mcm5p1f_cf_w_0_150_s_0_630=2.65e-11
.param mcm5p1f_ca_w_0_150_s_0_840=1.13e-04
.param mcm5p1f_cc_w_0_150_s_0_840=1.81e-11
.param mcm5p1f_cf_w_0_150_s_0_840=3.15e-11
.param mcm5p1f_ca_w_0_150_s_1_260=1.13e-04
.param mcm5p1f_cc_w_0_150_s_1_260=9.93e-12
.param mcm5p1f_cf_w_0_150_s_1_260=3.81e-11
.param mcm5p1f_ca_w_0_150_s_2_310=1.13e-04
.param mcm5p1f_cc_w_0_150_s_2_310=3.34e-12
.param mcm5p1f_cf_w_0_150_s_2_310=4.40e-11
.param mcm5p1f_ca_w_0_150_s_5_250=1.13e-04
.param mcm5p1f_cc_w_0_150_s_5_250=4.63e-13
.param mcm5p1f_cf_w_0_150_s_5_250=4.69e-11
.param mcm5p1f_ca_w_1_200_s_0_210=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_210=9.02e-11
.param mcm5p1f_cf_w_1_200_s_0_210=1.10e-11
.param mcm5p1f_ca_w_1_200_s_0_263=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_263=7.46e-11
.param mcm5p1f_cf_w_1_200_s_0_263=1.34e-11
.param mcm5p1f_ca_w_1_200_s_0_315=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_315=6.41e-11
.param mcm5p1f_cf_w_1_200_s_0_315=1.57e-11
.param mcm5p1f_ca_w_1_200_s_0_420=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_420=5.02e-11
.param mcm5p1f_cf_w_1_200_s_0_420=1.98e-11
.param mcm5p1f_ca_w_1_200_s_0_525=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_525=4.11e-11
.param mcm5p1f_cf_w_1_200_s_0_525=2.35e-11
.param mcm5p1f_ca_w_1_200_s_0_630=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_630=3.47e-11
.param mcm5p1f_cf_w_1_200_s_0_630=2.67e-11
.param mcm5p1f_ca_w_1_200_s_0_840=1.13e-04
.param mcm5p1f_cc_w_1_200_s_0_840=2.59e-11
.param mcm5p1f_cf_w_1_200_s_0_840=3.21e-11
.param mcm5p1f_ca_w_1_200_s_1_260=1.13e-04
.param mcm5p1f_cc_w_1_200_s_1_260=1.60e-11
.param mcm5p1f_cf_w_1_200_s_1_260=3.94e-11
.param mcm5p1f_ca_w_1_200_s_2_310=1.13e-04
.param mcm5p1f_cc_w_1_200_s_2_310=6.20e-12
.param mcm5p1f_cf_w_1_200_s_2_310=4.79e-11
.param mcm5p1f_ca_w_1_200_s_5_250=1.13e-04
.param mcm5p1f_cc_w_1_200_s_5_250=8.40e-13
.param mcm5p1f_cf_w_1_200_s_5_250=5.31e-11
.param mcrdlp1f_ca_w_0_150_s_0_210=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_210=7.57e-11
.param mcrdlp1f_cf_w_0_150_s_0_210=1.06e-11
.param mcrdlp1f_ca_w_0_150_s_0_263=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_263=6.15e-11
.param mcrdlp1f_cf_w_0_150_s_0_263=1.28e-11
.param mcrdlp1f_ca_w_0_150_s_0_315=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_315=5.24e-11
.param mcrdlp1f_cf_w_0_150_s_0_315=1.50e-11
.param mcrdlp1f_ca_w_0_150_s_0_420=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_420=3.98e-11
.param mcrdlp1f_cf_w_0_150_s_0_420=1.90e-11
.param mcrdlp1f_ca_w_0_150_s_0_525=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_525=3.23e-11
.param mcrdlp1f_cf_w_0_150_s_0_525=2.24e-11
.param mcrdlp1f_ca_w_0_150_s_0_630=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_630=2.69e-11
.param mcrdlp1f_cf_w_0_150_s_0_630=2.53e-11
.param mcrdlp1f_ca_w_0_150_s_0_840=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_0_840=1.95e-11
.param mcrdlp1f_cf_w_0_150_s_0_840=3.02e-11
.param mcrdlp1f_ca_w_0_150_s_1_260=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_1_260=1.11e-11
.param mcrdlp1f_cf_w_0_150_s_1_260=3.69e-11
.param mcrdlp1f_ca_w_0_150_s_2_310=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_2_310=4.42e-12
.param mcrdlp1f_cf_w_0_150_s_2_310=4.30e-11
.param mcrdlp1f_ca_w_0_150_s_5_250=1.09e-04
.param mcrdlp1f_cc_w_0_150_s_5_250=8.77e-13
.param mcrdlp1f_cf_w_0_150_s_5_250=4.65e-11
.param mcrdlp1f_ca_w_1_200_s_0_210=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_210=9.30e-11
.param mcrdlp1f_cf_w_1_200_s_0_210=1.05e-11
.param mcrdlp1f_ca_w_1_200_s_0_263=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_263=7.73e-11
.param mcrdlp1f_cf_w_1_200_s_0_263=1.28e-11
.param mcrdlp1f_ca_w_1_200_s_0_315=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_315=6.69e-11
.param mcrdlp1f_cf_w_1_200_s_0_315=1.50e-11
.param mcrdlp1f_ca_w_1_200_s_0_420=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_420=5.31e-11
.param mcrdlp1f_cf_w_1_200_s_0_420=1.90e-11
.param mcrdlp1f_ca_w_1_200_s_0_525=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_525=4.42e-11
.param mcrdlp1f_cf_w_1_200_s_0_525=2.25e-11
.param mcrdlp1f_ca_w_1_200_s_0_630=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_630=3.79e-11
.param mcrdlp1f_cf_w_1_200_s_0_630=2.56e-11
.param mcrdlp1f_ca_w_1_200_s_0_840=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_0_840=2.92e-11
.param mcrdlp1f_cf_w_1_200_s_0_840=3.08e-11
.param mcrdlp1f_ca_w_1_200_s_1_260=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_1_260=1.93e-11
.param mcrdlp1f_cf_w_1_200_s_1_260=3.80e-11
.param mcrdlp1f_ca_w_1_200_s_2_310=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_2_310=8.91e-12
.param mcrdlp1f_cf_w_1_200_s_2_310=4.71e-11
.param mcrdlp1f_ca_w_1_200_s_5_250=1.09e-04
.param mcrdlp1f_cc_w_1_200_s_5_250=2.15e-12
.param mcrdlp1f_cf_w_1_200_s_5_250=5.35e-11
.param mcm1l1f_ca_w_0_170_s_0_180=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_180=6.64e-11
.param mcm1l1f_cf_w_0_170_s_0_180=1.26e-11
.param mcm1l1f_ca_w_0_170_s_0_225=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_225=5.39e-11
.param mcm1l1f_cf_w_0_170_s_0_225=1.53e-11
.param mcm1l1f_ca_w_0_170_s_0_270=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_270=4.51e-11
.param mcm1l1f_cf_w_0_170_s_0_270=1.79e-11
.param mcm1l1f_ca_w_0_170_s_0_360=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_360=3.31e-11
.param mcm1l1f_cf_w_0_170_s_0_360=2.27e-11
.param mcm1l1f_ca_w_0_170_s_0_450=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_450=2.52e-11
.param mcm1l1f_cf_w_0_170_s_0_450=2.67e-11
.param mcm1l1f_ca_w_0_170_s_0_540=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_540=1.96e-11
.param mcm1l1f_cf_w_0_170_s_0_540=3.02e-11
.param mcm1l1f_ca_w_0_170_s_0_720=1.51e-04
.param mcm1l1f_cc_w_0_170_s_0_720=1.22e-11
.param mcm1l1f_cf_w_0_170_s_0_720=3.55e-11
.param mcm1l1f_ca_w_0_170_s_1_080=1.51e-04
.param mcm1l1f_cc_w_0_170_s_1_080=5.14e-12
.param mcm1l1f_cf_w_0_170_s_1_080=4.15e-11
.param mcm1l1f_ca_w_0_170_s_1_980=1.51e-04
.param mcm1l1f_cc_w_0_170_s_1_980=7.00e-13
.param mcm1l1f_cf_w_0_170_s_1_980=4.57e-11
.param mcm1l1f_ca_w_0_170_s_4_500=1.51e-04
.param mcm1l1f_cc_w_0_170_s_4_500=0.00e+00
.param mcm1l1f_cf_w_0_170_s_4_500=4.63e-11
.param mcm1l1f_ca_w_1_360_s_0_180=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_180=7.19e-11
.param mcm1l1f_cf_w_1_360_s_0_180=1.25e-11
.param mcm1l1f_ca_w_1_360_s_0_225=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_225=5.86e-11
.param mcm1l1f_cf_w_1_360_s_0_225=1.53e-11
.param mcm1l1f_ca_w_1_360_s_0_270=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_270=4.93e-11
.param mcm1l1f_cf_w_1_360_s_0_270=1.79e-11
.param mcm1l1f_ca_w_1_360_s_0_360=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_360=3.65e-11
.param mcm1l1f_cf_w_1_360_s_0_360=2.27e-11
.param mcm1l1f_ca_w_1_360_s_0_450=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_450=2.80e-11
.param mcm1l1f_cf_w_1_360_s_0_450=2.69e-11
.param mcm1l1f_ca_w_1_360_s_0_540=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_540=2.19e-11
.param mcm1l1f_cf_w_1_360_s_0_540=3.05e-11
.param mcm1l1f_ca_w_1_360_s_0_720=1.51e-04
.param mcm1l1f_cc_w_1_360_s_0_720=1.39e-11
.param mcm1l1f_cf_w_1_360_s_0_720=3.60e-11
.param mcm1l1f_ca_w_1_360_s_1_080=1.51e-04
.param mcm1l1f_cc_w_1_360_s_1_080=5.95e-12
.param mcm1l1f_cf_w_1_360_s_1_080=4.26e-11
.param mcm1l1f_ca_w_1_360_s_1_980=1.51e-04
.param mcm1l1f_cc_w_1_360_s_1_980=8.15e-13
.param mcm1l1f_cf_w_1_360_s_1_980=4.75e-11
.param mcm1l1f_ca_w_1_360_s_4_500=1.51e-04
.param mcm1l1f_cc_w_1_360_s_4_500=0.00e+00
.param mcm1l1f_cf_w_1_360_s_4_500=4.83e-11
.param mcm1l1d_ca_w_0_170_s_0_180=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_180=6.40e-11
.param mcm1l1d_cf_w_0_170_s_0_180=1.41e-11
.param mcm1l1d_ca_w_0_170_s_0_225=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_225=5.15e-11
.param mcm1l1d_cf_w_0_170_s_0_225=1.72e-11
.param mcm1l1d_ca_w_0_170_s_0_270=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_270=4.25e-11
.param mcm1l1d_cf_w_0_170_s_0_270=2.01e-11
.param mcm1l1d_ca_w_0_170_s_0_360=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_360=3.03e-11
.param mcm1l1d_cf_w_0_170_s_0_360=2.53e-11
.param mcm1l1d_ca_w_0_170_s_0_450=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_450=2.25e-11
.param mcm1l1d_cf_w_0_170_s_0_450=2.96e-11
.param mcm1l1d_ca_w_0_170_s_0_540=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_540=1.69e-11
.param mcm1l1d_cf_w_0_170_s_0_540=3.32e-11
.param mcm1l1d_ca_w_0_170_s_0_720=1.69e-04
.param mcm1l1d_cc_w_0_170_s_0_720=9.88e-12
.param mcm1l1d_cf_w_0_170_s_0_720=3.85e-11
.param mcm1l1d_ca_w_0_170_s_1_080=1.69e-04
.param mcm1l1d_cc_w_0_170_s_1_080=3.53e-12
.param mcm1l1d_cf_w_0_170_s_1_080=4.41e-11
.param mcm1l1d_ca_w_0_170_s_1_980=1.69e-04
.param mcm1l1d_cc_w_0_170_s_1_980=3.45e-13
.param mcm1l1d_cf_w_0_170_s_1_980=4.72e-11
.param mcm1l1d_ca_w_0_170_s_4_500=1.69e-04
.param mcm1l1d_cc_w_0_170_s_4_500=3.00e-14
.param mcm1l1d_cf_w_0_170_s_4_500=4.75e-11
.param mcm1l1d_ca_w_1_360_s_0_180=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_180=6.78e-11
.param mcm1l1d_cf_w_1_360_s_0_180=1.40e-11
.param mcm1l1d_ca_w_1_360_s_0_225=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_225=5.46e-11
.param mcm1l1d_cf_w_1_360_s_0_225=1.71e-11
.param mcm1l1d_ca_w_1_360_s_0_270=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_270=4.53e-11
.param mcm1l1d_cf_w_1_360_s_0_270=2.00e-11
.param mcm1l1d_ca_w_1_360_s_0_360=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_360=3.25e-11
.param mcm1l1d_cf_w_1_360_s_0_360=2.52e-11
.param mcm1l1d_ca_w_1_360_s_0_450=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_450=2.40e-11
.param mcm1l1d_cf_w_1_360_s_0_450=2.97e-11
.param mcm1l1d_ca_w_1_360_s_0_540=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_540=1.83e-11
.param mcm1l1d_cf_w_1_360_s_0_540=3.34e-11
.param mcm1l1d_ca_w_1_360_s_0_720=1.69e-04
.param mcm1l1d_cc_w_1_360_s_0_720=1.07e-11
.param mcm1l1d_cf_w_1_360_s_0_720=3.90e-11
.param mcm1l1d_ca_w_1_360_s_1_080=1.69e-04
.param mcm1l1d_cc_w_1_360_s_1_080=3.90e-12
.param mcm1l1d_cf_w_1_360_s_1_080=4.49e-11
.param mcm1l1d_ca_w_1_360_s_1_980=1.69e-04
.param mcm1l1d_cc_w_1_360_s_1_980=3.50e-13
.param mcm1l1d_cf_w_1_360_s_1_980=4.83e-11
.param mcm1l1d_ca_w_1_360_s_4_500=1.69e-04
.param mcm1l1d_cc_w_1_360_s_4_500=1.29e-26
.param mcm1l1d_cf_w_1_360_s_4_500=4.86e-11
.param mcm1l1p1_ca_w_0_170_s_0_180=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_180=5.98e-11
.param mcm1l1p1_cf_w_0_170_s_0_180=1.73e-11
.param mcm1l1p1_ca_w_0_170_s_0_225=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_225=4.72e-11
.param mcm1l1p1_cf_w_0_170_s_0_225=2.09e-11
.param mcm1l1p1_ca_w_0_170_s_0_270=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_270=3.81e-11
.param mcm1l1p1_cf_w_0_170_s_0_270=2.43e-11
.param mcm1l1p1_ca_w_0_170_s_0_360=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_360=2.60e-11
.param mcm1l1p1_cf_w_0_170_s_0_360=3.03e-11
.param mcm1l1p1_ca_w_0_170_s_0_450=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_450=1.82e-11
.param mcm1l1p1_cf_w_0_170_s_0_450=3.51e-11
.param mcm1l1p1_ca_w_0_170_s_0_540=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_540=1.30e-11
.param mcm1l1p1_cf_w_0_170_s_0_540=3.89e-11
.param mcm1l1p1_ca_w_0_170_s_0_720=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_0_720=6.77e-12
.param mcm1l1p1_cf_w_0_170_s_0_720=4.40e-11
.param mcm1l1p1_ca_w_0_170_s_1_080=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_1_080=1.87e-12
.param mcm1l1p1_cf_w_0_170_s_1_080=4.85e-11
.param mcm1l1p1_ca_w_0_170_s_1_980=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_1_980=9.50e-14
.param mcm1l1p1_cf_w_0_170_s_1_980=5.03e-11
.param mcm1l1p1_ca_w_0_170_s_4_500=2.08e-04
.param mcm1l1p1_cc_w_0_170_s_4_500=0.00e+00
.param mcm1l1p1_cf_w_0_170_s_4_500=5.04e-11
.param mcm1l1p1_ca_w_1_360_s_0_180=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_180=6.16e-11
.param mcm1l1p1_cf_w_1_360_s_0_180=1.71e-11
.param mcm1l1p1_ca_w_1_360_s_0_225=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_225=4.86e-11
.param mcm1l1p1_cf_w_1_360_s_0_225=2.08e-11
.param mcm1l1p1_ca_w_1_360_s_0_270=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_270=3.93e-11
.param mcm1l1p1_cf_w_1_360_s_0_270=2.43e-11
.param mcm1l1p1_ca_w_1_360_s_0_360=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_360=2.69e-11
.param mcm1l1p1_cf_w_1_360_s_0_360=3.02e-11
.param mcm1l1p1_ca_w_1_360_s_0_450=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_450=1.88e-11
.param mcm1l1p1_cf_w_1_360_s_0_450=3.52e-11
.param mcm1l1p1_ca_w_1_360_s_0_540=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_540=1.35e-11
.param mcm1l1p1_cf_w_1_360_s_0_540=3.90e-11
.param mcm1l1p1_ca_w_1_360_s_0_720=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_0_720=7.00e-12
.param mcm1l1p1_cf_w_1_360_s_0_720=4.43e-11
.param mcm1l1p1_ca_w_1_360_s_1_080=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_1_080=1.95e-12
.param mcm1l1p1_cf_w_1_360_s_1_080=4.90e-11
.param mcm1l1p1_ca_w_1_360_s_1_980=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_1_980=1.50e-13
.param mcm1l1p1_cf_w_1_360_s_1_980=5.08e-11
.param mcm1l1p1_ca_w_1_360_s_4_500=2.08e-04
.param mcm1l1p1_cc_w_1_360_s_4_500=0.00e+00
.param mcm1l1p1_cf_w_1_360_s_4_500=5.08e-11
.param mcm2l1f_ca_w_0_170_s_0_180=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_180=7.49e-11
.param mcm2l1f_cf_w_0_170_s_0_180=6.47e-12
.param mcm2l1f_ca_w_0_170_s_0_225=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_225=6.27e-11
.param mcm2l1f_cf_w_0_170_s_0_225=8.02e-12
.param mcm2l1f_ca_w_0_170_s_0_270=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_270=5.41e-11
.param mcm2l1f_cf_w_0_170_s_0_270=9.48e-12
.param mcm2l1f_ca_w_0_170_s_0_360=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_360=4.24e-11
.param mcm2l1f_cf_w_0_170_s_0_360=1.24e-11
.param mcm2l1f_ca_w_0_170_s_0_450=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_450=3.45e-11
.param mcm2l1f_cf_w_0_170_s_0_450=1.50e-11
.param mcm2l1f_ca_w_0_170_s_0_540=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_540=2.87e-11
.param mcm2l1f_cf_w_0_170_s_0_540=1.75e-11
.param mcm2l1f_ca_w_0_170_s_0_720=7.40e-05
.param mcm2l1f_cc_w_0_170_s_0_720=2.06e-11
.param mcm2l1f_cf_w_0_170_s_0_720=2.17e-11
.param mcm2l1f_ca_w_0_170_s_1_080=7.40e-05
.param mcm2l1f_cc_w_0_170_s_1_080=1.13e-11
.param mcm2l1f_cf_w_0_170_s_1_080=2.79e-11
.param mcm2l1f_ca_w_0_170_s_1_980=7.40e-05
.param mcm2l1f_cc_w_0_170_s_1_980=2.81e-12
.param mcm2l1f_cf_w_0_170_s_1_980=3.50e-11
.param mcm2l1f_ca_w_0_170_s_4_500=7.40e-05
.param mcm2l1f_cc_w_0_170_s_4_500=9.50e-14
.param mcm2l1f_cf_w_0_170_s_4_500=3.76e-11
.param mcm2l1f_ca_w_1_360_s_0_180=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_180=8.41e-11
.param mcm2l1f_cf_w_1_360_s_0_180=6.43e-12
.param mcm2l1f_ca_w_1_360_s_0_225=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_225=7.09e-11
.param mcm2l1f_cf_w_1_360_s_0_225=7.97e-12
.param mcm2l1f_ca_w_1_360_s_0_270=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_270=6.14e-11
.param mcm2l1f_cf_w_1_360_s_0_270=9.48e-12
.param mcm2l1f_ca_w_1_360_s_0_360=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_360=4.83e-11
.param mcm2l1f_cf_w_1_360_s_0_360=1.24e-11
.param mcm2l1f_ca_w_1_360_s_0_450=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_450=3.94e-11
.param mcm2l1f_cf_w_1_360_s_0_450=1.51e-11
.param mcm2l1f_ca_w_1_360_s_0_540=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_540=3.29e-11
.param mcm2l1f_cf_w_1_360_s_0_540=1.76e-11
.param mcm2l1f_ca_w_1_360_s_0_720=7.40e-05
.param mcm2l1f_cc_w_1_360_s_0_720=2.37e-11
.param mcm2l1f_cf_w_1_360_s_0_720=2.21e-11
.param mcm2l1f_ca_w_1_360_s_1_080=7.40e-05
.param mcm2l1f_cc_w_1_360_s_1_080=1.32e-11
.param mcm2l1f_cf_w_1_360_s_1_080=2.88e-11
.param mcm2l1f_ca_w_1_360_s_1_980=7.40e-05
.param mcm2l1f_cc_w_1_360_s_1_980=3.32e-12
.param mcm2l1f_cf_w_1_360_s_1_980=3.70e-11
.param mcm2l1f_ca_w_1_360_s_4_500=7.40e-05
.param mcm2l1f_cc_w_1_360_s_4_500=1.30e-13
.param mcm2l1f_cf_w_1_360_s_4_500=4.01e-11
.param mcm2l1d_ca_w_0_170_s_0_180=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_180=7.24e-11
.param mcm2l1d_cf_w_0_170_s_0_180=8.03e-12
.param mcm2l1d_ca_w_0_170_s_0_225=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_225=6.02e-11
.param mcm2l1d_cf_w_0_170_s_0_225=9.90e-12
.param mcm2l1d_ca_w_0_170_s_0_270=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_270=5.14e-11
.param mcm2l1d_cf_w_0_170_s_0_270=1.17e-11
.param mcm2l1d_ca_w_0_170_s_0_360=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_360=3.94e-11
.param mcm2l1d_cf_w_0_170_s_0_360=1.52e-11
.param mcm2l1d_ca_w_0_170_s_0_450=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_450=3.15e-11
.param mcm2l1d_cf_w_0_170_s_0_450=1.83e-11
.param mcm2l1d_ca_w_0_170_s_0_540=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_540=2.56e-11
.param mcm2l1d_cf_w_0_170_s_0_540=2.11e-11
.param mcm2l1d_ca_w_0_170_s_0_720=9.23e-05
.param mcm2l1d_cc_w_0_170_s_0_720=1.76e-11
.param mcm2l1d_cf_w_0_170_s_0_720=2.58e-11
.param mcm2l1d_ca_w_0_170_s_1_080=9.23e-05
.param mcm2l1d_cc_w_0_170_s_1_080=8.77e-12
.param mcm2l1d_cf_w_0_170_s_1_080=3.23e-11
.param mcm2l1d_ca_w_0_170_s_1_980=9.23e-05
.param mcm2l1d_cc_w_0_170_s_1_980=1.71e-12
.param mcm2l1d_cf_w_0_170_s_1_980=3.85e-11
.param mcm2l1d_ca_w_0_170_s_4_500=9.23e-05
.param mcm2l1d_cc_w_0_170_s_4_500=4.50e-14
.param mcm2l1d_cf_w_0_170_s_4_500=4.01e-11
.param mcm2l1d_ca_w_1_360_s_0_180=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_180=7.96e-11
.param mcm2l1d_cf_w_1_360_s_0_180=7.99e-12
.param mcm2l1d_ca_w_1_360_s_0_225=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_225=6.65e-11
.param mcm2l1d_cf_w_1_360_s_0_225=9.88e-12
.param mcm2l1d_ca_w_1_360_s_0_270=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_270=5.70e-11
.param mcm2l1d_cf_w_1_360_s_0_270=1.17e-11
.param mcm2l1d_ca_w_1_360_s_0_360=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_360=4.39e-11
.param mcm2l1d_cf_w_1_360_s_0_360=1.52e-11
.param mcm2l1d_ca_w_1_360_s_0_450=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_450=3.51e-11
.param mcm2l1d_cf_w_1_360_s_0_450=1.84e-11
.param mcm2l1d_ca_w_1_360_s_0_540=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_540=2.87e-11
.param mcm2l1d_cf_w_1_360_s_0_540=2.13e-11
.param mcm2l1d_ca_w_1_360_s_0_720=9.23e-05
.param mcm2l1d_cc_w_1_360_s_0_720=1.98e-11
.param mcm2l1d_cf_w_1_360_s_0_720=2.63e-11
.param mcm2l1d_ca_w_1_360_s_1_080=9.23e-05
.param mcm2l1d_cc_w_1_360_s_1_080=1.01e-11
.param mcm2l1d_cf_w_1_360_s_1_080=3.33e-11
.param mcm2l1d_ca_w_1_360_s_1_980=9.23e-05
.param mcm2l1d_cc_w_1_360_s_1_980=1.97e-12
.param mcm2l1d_cf_w_1_360_s_1_980=4.04e-11
.param mcm2l1d_ca_w_1_360_s_4_500=9.23e-05
.param mcm2l1d_cc_w_1_360_s_4_500=9.50e-14
.param mcm2l1d_cf_w_1_360_s_4_500=4.23e-11
.param mcm2l1p1_ca_w_0_170_s_0_180=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_180=6.82e-11
.param mcm2l1p1_cf_w_0_170_s_0_180=1.12e-11
.param mcm2l1p1_ca_w_0_170_s_0_225=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_225=5.56e-11
.param mcm2l1p1_cf_w_0_170_s_0_225=1.38e-11
.param mcm2l1p1_ca_w_0_170_s_0_270=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_270=4.68e-11
.param mcm2l1p1_cf_w_0_170_s_0_270=1.62e-11
.param mcm2l1p1_ca_w_0_170_s_0_360=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_360=3.47e-11
.param mcm2l1p1_cf_w_0_170_s_0_360=2.08e-11
.param mcm2l1p1_ca_w_0_170_s_0_450=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_450=2.68e-11
.param mcm2l1p1_cf_w_0_170_s_0_450=2.46e-11
.param mcm2l1p1_ca_w_0_170_s_0_540=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_540=2.10e-11
.param mcm2l1p1_cf_w_0_170_s_0_540=2.80e-11
.param mcm2l1p1_ca_w_0_170_s_0_720=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_0_720=1.34e-11
.param mcm2l1p1_cf_w_0_170_s_0_720=3.33e-11
.param mcm2l1p1_ca_w_0_170_s_1_080=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_1_080=5.79e-12
.param mcm2l1p1_cf_w_0_170_s_1_080=3.95e-11
.param mcm2l1p1_ca_w_0_170_s_1_980=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_1_980=8.00e-13
.param mcm2l1p1_cf_w_0_170_s_1_980=4.41e-11
.param mcm2l1p1_ca_w_0_170_s_4_500=1.31e-04
.param mcm2l1p1_cc_w_0_170_s_4_500=5.00e-15
.param mcm2l1p1_cf_w_0_170_s_4_500=4.49e-11
.param mcm2l1p1_ca_w_1_360_s_0_180=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_180=7.38e-11
.param mcm2l1p1_cf_w_1_360_s_0_180=1.12e-11
.param mcm2l1p1_ca_w_1_360_s_0_225=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_225=6.07e-11
.param mcm2l1p1_cf_w_1_360_s_0_225=1.37e-11
.param mcm2l1p1_ca_w_1_360_s_0_270=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_270=5.13e-11
.param mcm2l1p1_cf_w_1_360_s_0_270=1.62e-11
.param mcm2l1p1_ca_w_1_360_s_0_360=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_360=3.83e-11
.param mcm2l1p1_cf_w_1_360_s_0_360=2.07e-11
.param mcm2l1p1_ca_w_1_360_s_0_450=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_450=2.97e-11
.param mcm2l1p1_cf_w_1_360_s_0_450=2.47e-11
.param mcm2l1p1_ca_w_1_360_s_0_540=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_540=2.35e-11
.param mcm2l1p1_cf_w_1_360_s_0_540=2.82e-11
.param mcm2l1p1_ca_w_1_360_s_0_720=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_0_720=1.52e-11
.param mcm2l1p1_cf_w_1_360_s_0_720=3.37e-11
.param mcm2l1p1_ca_w_1_360_s_1_080=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_1_080=6.72e-12
.param mcm2l1p1_cf_w_1_360_s_1_080=4.06e-11
.param mcm2l1p1_ca_w_1_360_s_1_980=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_1_980=9.95e-13
.param mcm2l1p1_cf_w_1_360_s_1_980=4.59e-11
.param mcm2l1p1_ca_w_1_360_s_4_500=1.31e-04
.param mcm2l1p1_cc_w_1_360_s_4_500=6.00e-14
.param mcm2l1p1_cf_w_1_360_s_4_500=4.69e-11
.param mcm3l1f_ca_w_0_170_s_0_180=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_180=7.71e-11
.param mcm3l1f_cf_w_0_170_s_0_180=5.03e-12
.param mcm3l1f_ca_w_0_170_s_0_225=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_225=6.52e-11
.param mcm3l1f_cf_w_0_170_s_0_225=6.25e-12
.param mcm3l1f_ca_w_0_170_s_0_270=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_270=5.70e-11
.param mcm3l1f_cf_w_0_170_s_0_270=7.41e-12
.param mcm3l1f_ca_w_0_170_s_0_360=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_360=4.55e-11
.param mcm3l1f_cf_w_0_170_s_0_360=9.84e-12
.param mcm3l1f_ca_w_0_170_s_0_450=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_450=3.81e-11
.param mcm3l1f_cf_w_0_170_s_0_450=1.18e-11
.param mcm3l1f_ca_w_0_170_s_0_540=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_540=3.22e-11
.param mcm3l1f_cf_w_0_170_s_0_540=1.40e-11
.param mcm3l1f_ca_w_0_170_s_0_720=5.71e-05
.param mcm3l1f_cc_w_0_170_s_0_720=2.43e-11
.param mcm3l1f_cf_w_0_170_s_0_720=1.76e-11
.param mcm3l1f_ca_w_0_170_s_1_080=5.71e-05
.param mcm3l1f_cc_w_0_170_s_1_080=1.48e-11
.param mcm3l1f_cf_w_0_170_s_1_080=2.32e-11
.param mcm3l1f_ca_w_0_170_s_1_980=5.71e-05
.param mcm3l1f_cc_w_0_170_s_1_980=4.96e-12
.param mcm3l1f_cf_w_0_170_s_1_980=3.10e-11
.param mcm3l1f_ca_w_0_170_s_4_500=5.71e-05
.param mcm3l1f_cc_w_0_170_s_4_500=3.10e-13
.param mcm3l1f_cf_w_0_170_s_4_500=3.53e-11
.param mcm3l1f_ca_w_1_360_s_0_180=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_180=9.02e-11
.param mcm3l1f_cf_w_1_360_s_0_180=5.01e-12
.param mcm3l1f_ca_w_1_360_s_0_225=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_225=7.69e-11
.param mcm3l1f_cf_w_1_360_s_0_225=6.22e-12
.param mcm3l1f_ca_w_1_360_s_0_270=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_270=6.75e-11
.param mcm3l1f_cf_w_1_360_s_0_270=7.41e-12
.param mcm3l1f_ca_w_1_360_s_0_360=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_360=5.44e-11
.param mcm3l1f_cf_w_1_360_s_0_360=9.72e-12
.param mcm3l1f_ca_w_1_360_s_0_450=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_450=4.55e-11
.param mcm3l1f_cf_w_1_360_s_0_450=1.19e-11
.param mcm3l1f_ca_w_1_360_s_0_540=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_540=3.89e-11
.param mcm3l1f_cf_w_1_360_s_0_540=1.40e-11
.param mcm3l1f_ca_w_1_360_s_0_720=5.71e-05
.param mcm3l1f_cc_w_1_360_s_0_720=2.95e-11
.param mcm3l1f_cf_w_1_360_s_0_720=1.78e-11
.param mcm3l1f_ca_w_1_360_s_1_080=5.71e-05
.param mcm3l1f_cc_w_1_360_s_1_080=1.83e-11
.param mcm3l1f_cf_w_1_360_s_1_080=2.40e-11
.param mcm3l1f_ca_w_1_360_s_1_980=5.71e-05
.param mcm3l1f_cc_w_1_360_s_1_980=6.38e-12
.param mcm3l1f_cf_w_1_360_s_1_980=3.31e-11
.param mcm3l1f_ca_w_1_360_s_4_500=5.71e-05
.param mcm3l1f_cc_w_1_360_s_4_500=3.95e-13
.param mcm3l1f_cf_w_1_360_s_4_500=3.86e-11
.param mcm3l1d_ca_w_0_170_s_0_180=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_180=7.47e-11
.param mcm3l1d_cf_w_0_170_s_0_180=6.60e-12
.param mcm3l1d_ca_w_0_170_s_0_225=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_225=6.26e-11
.param mcm3l1d_cf_w_0_170_s_0_225=8.16e-12
.param mcm3l1d_ca_w_0_170_s_0_270=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_270=5.43e-11
.param mcm3l1d_cf_w_0_170_s_0_270=9.66e-12
.param mcm3l1d_ca_w_0_170_s_0_360=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_360=4.25e-11
.param mcm3l1d_cf_w_0_170_s_0_360=1.27e-11
.param mcm3l1d_ca_w_0_170_s_0_450=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_450=3.49e-11
.param mcm3l1d_cf_w_0_170_s_0_450=1.52e-11
.param mcm3l1d_ca_w_0_170_s_0_540=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_540=2.90e-11
.param mcm3l1d_cf_w_0_170_s_0_540=1.78e-11
.param mcm3l1d_ca_w_0_170_s_0_720=7.54e-05
.param mcm3l1d_cc_w_0_170_s_0_720=2.10e-11
.param mcm3l1d_cf_w_0_170_s_0_720=2.20e-11
.param mcm3l1d_ca_w_0_170_s_1_080=7.54e-05
.param mcm3l1d_cc_w_0_170_s_1_080=1.19e-11
.param mcm3l1d_cf_w_0_170_s_1_080=2.82e-11
.param mcm3l1d_ca_w_0_170_s_1_980=7.54e-05
.param mcm3l1d_cc_w_0_170_s_1_980=3.34e-12
.param mcm3l1d_cf_w_0_170_s_1_980=3.54e-11
.param mcm3l1d_ca_w_0_170_s_4_500=7.54e-05
.param mcm3l1d_cc_w_0_170_s_4_500=1.60e-13
.param mcm3l1d_cf_w_0_170_s_4_500=3.85e-11
.param mcm3l1d_ca_w_1_360_s_0_180=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_180=8.58e-11
.param mcm3l1d_cf_w_1_360_s_0_180=6.57e-12
.param mcm3l1d_ca_w_1_360_s_0_225=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_225=7.25e-11
.param mcm3l1d_cf_w_1_360_s_0_225=8.14e-12
.param mcm3l1d_ca_w_1_360_s_0_270=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_270=6.31e-11
.param mcm3l1d_cf_w_1_360_s_0_270=9.67e-12
.param mcm3l1d_ca_w_1_360_s_0_360=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_360=5.01e-11
.param mcm3l1d_cf_w_1_360_s_0_360=1.26e-11
.param mcm3l1d_ca_w_1_360_s_0_450=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_450=4.12e-11
.param mcm3l1d_cf_w_1_360_s_0_450=1.53e-11
.param mcm3l1d_ca_w_1_360_s_0_540=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_540=3.46e-11
.param mcm3l1d_cf_w_1_360_s_0_540=1.79e-11
.param mcm3l1d_ca_w_1_360_s_0_720=7.54e-05
.param mcm3l1d_cc_w_1_360_s_0_720=2.55e-11
.param mcm3l1d_cf_w_1_360_s_0_720=2.24e-11
.param mcm3l1d_ca_w_1_360_s_1_080=7.54e-05
.param mcm3l1d_cc_w_1_360_s_1_080=1.48e-11
.param mcm3l1d_cf_w_1_360_s_1_080=2.92e-11
.param mcm3l1d_ca_w_1_360_s_1_980=7.54e-05
.param mcm3l1d_cc_w_1_360_s_1_980=4.42e-12
.param mcm3l1d_cf_w_1_360_s_1_980=3.78e-11
.param mcm3l1d_ca_w_1_360_s_4_500=7.54e-05
.param mcm3l1d_cc_w_1_360_s_4_500=1.80e-13
.param mcm3l1d_cf_w_1_360_s_4_500=4.19e-11
.param mcm3l1p1_ca_w_0_170_s_0_180=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_180=7.05e-11
.param mcm3l1p1_cf_w_0_170_s_0_180=9.84e-12
.param mcm3l1p1_ca_w_0_170_s_0_225=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_225=5.82e-11
.param mcm3l1p1_cf_w_0_170_s_0_225=1.21e-11
.param mcm3l1p1_ca_w_0_170_s_0_270=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_270=4.96e-11
.param mcm3l1p1_cf_w_0_170_s_0_270=1.42e-11
.param mcm3l1p1_ca_w_0_170_s_0_360=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_360=3.76e-11
.param mcm3l1p1_cf_w_0_170_s_0_360=1.84e-11
.param mcm3l1p1_ca_w_0_170_s_0_450=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_450=3.00e-11
.param mcm3l1p1_cf_w_0_170_s_0_450=2.18e-11
.param mcm3l1p1_ca_w_0_170_s_0_540=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_540=2.42e-11
.param mcm3l1p1_cf_w_0_170_s_0_540=2.51e-11
.param mcm3l1p1_ca_w_0_170_s_0_720=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_0_720=1.64e-11
.param mcm3l1p1_cf_w_0_170_s_0_720=3.01e-11
.param mcm3l1p1_ca_w_0_170_s_1_080=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_1_080=8.31e-12
.param mcm3l1p1_cf_w_0_170_s_1_080=3.65e-11
.param mcm3l1p1_ca_w_0_170_s_1_980=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_1_980=1.89e-12
.param mcm3l1p1_cf_w_0_170_s_1_980=4.22e-11
.param mcm3l1p1_ca_w_0_170_s_4_500=1.14e-04
.param mcm3l1p1_cc_w_0_170_s_4_500=7.00e-14
.param mcm3l1p1_cf_w_0_170_s_4_500=4.40e-11
.param mcm3l1p1_ca_w_1_360_s_0_180=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_180=7.98e-11
.param mcm3l1p1_cf_w_1_360_s_0_180=9.83e-12
.param mcm3l1p1_ca_w_1_360_s_0_225=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_225=6.68e-11
.param mcm3l1p1_cf_w_1_360_s_0_225=1.21e-11
.param mcm3l1p1_ca_w_1_360_s_0_270=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_270=5.72e-11
.param mcm3l1p1_cf_w_1_360_s_0_270=1.42e-11
.param mcm3l1p1_ca_w_1_360_s_0_360=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_360=4.43e-11
.param mcm3l1p1_cf_w_1_360_s_0_360=1.83e-11
.param mcm3l1p1_ca_w_1_360_s_0_450=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_450=3.56e-11
.param mcm3l1p1_cf_w_1_360_s_0_450=2.19e-11
.param mcm3l1p1_ca_w_1_360_s_0_540=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_540=2.92e-11
.param mcm3l1p1_cf_w_1_360_s_0_540=2.52e-11
.param mcm3l1p1_ca_w_1_360_s_0_720=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_0_720=2.05e-11
.param mcm3l1p1_cf_w_1_360_s_0_720=3.05e-11
.param mcm3l1p1_ca_w_1_360_s_1_080=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_1_080=1.09e-11
.param mcm3l1p1_cf_w_1_360_s_1_080=3.78e-11
.param mcm3l1p1_ca_w_1_360_s_1_980=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_1_980=2.72e-12
.param mcm3l1p1_cf_w_1_360_s_1_980=4.51e-11
.param mcm3l1p1_ca_w_1_360_s_4_500=1.14e-04
.param mcm3l1p1_cc_w_1_360_s_4_500=1.05e-13
.param mcm3l1p1_cf_w_1_360_s_4_500=4.77e-11
.param mcm4l1f_ca_w_0_170_s_0_180=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_180=7.83e-11
.param mcm4l1f_cf_w_0_170_s_0_180=4.30e-12
.param mcm4l1f_ca_w_0_170_s_0_225=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_225=6.66e-11
.param mcm4l1f_cf_w_0_170_s_0_225=5.34e-12
.param mcm4l1f_ca_w_0_170_s_0_270=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_270=5.85e-11
.param mcm4l1f_cf_w_0_170_s_0_270=6.33e-12
.param mcm4l1f_ca_w_0_170_s_0_360=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_360=4.72e-11
.param mcm4l1f_cf_w_0_170_s_0_360=8.48e-12
.param mcm4l1f_ca_w_0_170_s_0_450=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_450=4.00e-11
.param mcm4l1f_cf_w_0_170_s_0_450=1.02e-11
.param mcm4l1f_ca_w_0_170_s_0_540=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_540=3.43e-11
.param mcm4l1f_cf_w_0_170_s_0_540=1.21e-11
.param mcm4l1f_ca_w_0_170_s_0_720=4.86e-05
.param mcm4l1f_cc_w_0_170_s_0_720=2.66e-11
.param mcm4l1f_cf_w_0_170_s_0_720=1.54e-11
.param mcm4l1f_ca_w_0_170_s_1_080=4.86e-05
.param mcm4l1f_cc_w_0_170_s_1_080=1.73e-11
.param mcm4l1f_cf_w_0_170_s_1_080=2.06e-11
.param mcm4l1f_ca_w_0_170_s_1_980=4.86e-05
.param mcm4l1f_cc_w_0_170_s_1_980=6.95e-12
.param mcm4l1f_cf_w_0_170_s_1_980=2.83e-11
.param mcm4l1f_ca_w_0_170_s_4_500=4.86e-05
.param mcm4l1f_cc_w_0_170_s_4_500=8.15e-13
.param mcm4l1f_cf_w_0_170_s_4_500=3.39e-11
.param mcm4l1f_ca_w_1_360_s_0_180=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_180=9.45e-11
.param mcm4l1f_cf_w_1_360_s_0_180=4.29e-12
.param mcm4l1f_ca_w_1_360_s_0_225=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_225=8.12e-11
.param mcm4l1f_cf_w_1_360_s_0_225=5.32e-12
.param mcm4l1f_ca_w_1_360_s_0_270=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_270=7.19e-11
.param mcm4l1f_cf_w_1_360_s_0_270=6.35e-12
.param mcm4l1f_ca_w_1_360_s_0_360=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_360=5.89e-11
.param mcm4l1f_cf_w_1_360_s_0_360=8.33e-12
.param mcm4l1f_ca_w_1_360_s_0_450=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_450=5.00e-11
.param mcm4l1f_cf_w_1_360_s_0_450=1.02e-11
.param mcm4l1f_ca_w_1_360_s_0_540=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_540=4.35e-11
.param mcm4l1f_cf_w_1_360_s_0_540=1.21e-11
.param mcm4l1f_ca_w_1_360_s_0_720=4.86e-05
.param mcm4l1f_cc_w_1_360_s_0_720=3.41e-11
.param mcm4l1f_cf_w_1_360_s_0_720=1.54e-11
.param mcm4l1f_ca_w_1_360_s_1_080=4.86e-05
.param mcm4l1f_cc_w_1_360_s_1_080=2.28e-11
.param mcm4l1f_cf_w_1_360_s_1_080=2.11e-11
.param mcm4l1f_ca_w_1_360_s_1_980=4.86e-05
.param mcm4l1f_cc_w_1_360_s_1_980=9.76e-12
.param mcm4l1f_cf_w_1_360_s_1_980=3.03e-11
.param mcm4l1f_ca_w_1_360_s_4_500=4.86e-05
.param mcm4l1f_cc_w_1_360_s_4_500=1.23e-12
.param mcm4l1f_cf_w_1_360_s_4_500=3.80e-11
.param mcm4l1d_ca_w_0_170_s_0_180=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_180=7.59e-11
.param mcm4l1d_cf_w_0_170_s_0_180=5.86e-12
.param mcm4l1d_ca_w_0_170_s_0_225=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_225=6.39e-11
.param mcm4l1d_cf_w_0_170_s_0_225=7.26e-12
.param mcm4l1d_ca_w_0_170_s_0_270=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_270=5.58e-11
.param mcm4l1d_cf_w_0_170_s_0_270=8.60e-12
.param mcm4l1d_ca_w_0_170_s_0_360=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_360=4.42e-11
.param mcm4l1d_cf_w_0_170_s_0_360=1.14e-11
.param mcm4l1d_ca_w_0_170_s_0_450=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_450=3.68e-11
.param mcm4l1d_cf_w_0_170_s_0_450=1.36e-11
.param mcm4l1d_ca_w_0_170_s_0_540=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_540=3.09e-11
.param mcm4l1d_cf_w_0_170_s_0_540=1.61e-11
.param mcm4l1d_ca_w_0_170_s_0_720=6.70e-05
.param mcm4l1d_cc_w_0_170_s_0_720=2.31e-11
.param mcm4l1d_cf_w_0_170_s_0_720=2.00e-11
.param mcm4l1d_ca_w_0_170_s_1_080=6.70e-05
.param mcm4l1d_cc_w_0_170_s_1_080=1.40e-11
.param mcm4l1d_cf_w_0_170_s_1_080=2.60e-11
.param mcm4l1d_ca_w_0_170_s_1_980=6.70e-05
.param mcm4l1d_cc_w_0_170_s_1_980=4.91e-12
.param mcm4l1d_cf_w_0_170_s_1_980=3.35e-11
.param mcm4l1d_ca_w_0_170_s_4_500=6.70e-05
.param mcm4l1d_cc_w_0_170_s_4_500=4.70e-13
.param mcm4l1d_cf_w_0_170_s_4_500=3.76e-11
.param mcm4l1d_ca_w_1_360_s_0_180=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_180=9.01e-11
.param mcm4l1d_cf_w_1_360_s_0_180=5.85e-12
.param mcm4l1d_ca_w_1_360_s_0_225=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_225=7.69e-11
.param mcm4l1d_cf_w_1_360_s_0_225=7.25e-12
.param mcm4l1d_ca_w_1_360_s_0_270=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_270=6.75e-11
.param mcm4l1d_cf_w_1_360_s_0_270=8.62e-12
.param mcm4l1d_ca_w_1_360_s_0_360=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_360=5.45e-11
.param mcm4l1d_cf_w_1_360_s_0_360=1.12e-11
.param mcm4l1d_ca_w_1_360_s_0_450=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_450=4.57e-11
.param mcm4l1d_cf_w_1_360_s_0_450=1.37e-11
.param mcm4l1d_ca_w_1_360_s_0_540=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_540=3.92e-11
.param mcm4l1d_cf_w_1_360_s_0_540=1.61e-11
.param mcm4l1d_ca_w_1_360_s_0_720=6.70e-05
.param mcm4l1d_cc_w_1_360_s_0_720=2.99e-11
.param mcm4l1d_cf_w_1_360_s_0_720=2.02e-11
.param mcm4l1d_ca_w_1_360_s_1_080=6.70e-05
.param mcm4l1d_cc_w_1_360_s_1_080=1.90e-11
.param mcm4l1d_cf_w_1_360_s_1_080=2.68e-11
.param mcm4l1d_ca_w_1_360_s_1_980=6.70e-05
.param mcm4l1d_cc_w_1_360_s_1_980=7.34e-12
.param mcm4l1d_cf_w_1_360_s_1_980=3.60e-11
.param mcm4l1d_ca_w_1_360_s_4_500=6.70e-05
.param mcm4l1d_cc_w_1_360_s_4_500=7.80e-13
.param mcm4l1d_cf_w_1_360_s_4_500=4.22e-11
.param mcm4l1p1_ca_w_0_170_s_0_180=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_180=7.17e-11
.param mcm4l1p1_cf_w_0_170_s_0_180=9.12e-12
.param mcm4l1p1_ca_w_0_170_s_0_225=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_225=5.95e-11
.param mcm4l1p1_cf_w_0_170_s_0_225=1.12e-11
.param mcm4l1p1_ca_w_0_170_s_0_270=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_270=5.11e-11
.param mcm4l1p1_cf_w_0_170_s_0_270=1.32e-11
.param mcm4l1p1_ca_w_0_170_s_0_360=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_360=3.92e-11
.param mcm4l1p1_cf_w_0_170_s_0_360=1.72e-11
.param mcm4l1p1_ca_w_0_170_s_0_450=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_450=3.18e-11
.param mcm4l1p1_cf_w_0_170_s_0_450=2.03e-11
.param mcm4l1p1_ca_w_0_170_s_0_540=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_540=2.59e-11
.param mcm4l1p1_cf_w_0_170_s_0_540=2.35e-11
.param mcm4l1p1_ca_w_0_170_s_0_720=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_0_720=1.83e-11
.param mcm4l1p1_cf_w_0_170_s_0_720=2.83e-11
.param mcm4l1p1_ca_w_0_170_s_1_080=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_1_080=1.00e-11
.param mcm4l1p1_cf_w_0_170_s_1_080=3.48e-11
.param mcm4l1p1_ca_w_0_170_s_1_980=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_1_980=2.96e-12
.param mcm4l1p1_cf_w_0_170_s_1_980=4.10e-11
.param mcm4l1p1_ca_w_0_170_s_4_500=1.06e-04
.param mcm4l1p1_cc_w_0_170_s_4_500=2.65e-13
.param mcm4l1p1_cf_w_0_170_s_4_500=4.37e-11
.param mcm4l1p1_ca_w_1_360_s_0_180=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_180=8.41e-11
.param mcm4l1p1_cf_w_1_360_s_0_180=9.16e-12
.param mcm4l1p1_ca_w_1_360_s_0_225=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_225=7.11e-11
.param mcm4l1p1_cf_w_1_360_s_0_225=1.13e-11
.param mcm4l1p1_ca_w_1_360_s_0_270=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_270=6.17e-11
.param mcm4l1p1_cf_w_1_360_s_0_270=1.33e-11
.param mcm4l1p1_ca_w_1_360_s_0_360=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_360=4.88e-11
.param mcm4l1p1_cf_w_1_360_s_0_360=1.70e-11
.param mcm4l1p1_ca_w_1_360_s_0_450=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_450=4.00e-11
.param mcm4l1p1_cf_w_1_360_s_0_450=2.05e-11
.param mcm4l1p1_ca_w_1_360_s_0_540=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_540=3.37e-11
.param mcm4l1p1_cf_w_1_360_s_0_540=2.36e-11
.param mcm4l1p1_ca_w_1_360_s_0_720=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_0_720=2.48e-11
.param mcm4l1p1_cf_w_1_360_s_0_720=2.87e-11
.param mcm4l1p1_ca_w_1_360_s_1_080=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_1_080=1.48e-11
.param mcm4l1p1_cf_w_1_360_s_1_080=3.61e-11
.param mcm4l1p1_ca_w_1_360_s_1_980=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_1_980=5.02e-12
.param mcm4l1p1_cf_w_1_360_s_1_980=4.46e-11
.param mcm4l1p1_ca_w_1_360_s_4_500=1.06e-04
.param mcm4l1p1_cc_w_1_360_s_4_500=4.55e-13
.param mcm4l1p1_cf_w_1_360_s_4_500=4.90e-11
.param mcm5l1f_ca_w_0_170_s_0_180=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_180=7.88e-11
.param mcm5l1f_cf_w_0_170_s_0_180=3.98e-12
.param mcm5l1f_ca_w_0_170_s_0_225=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_225=6.71e-11
.param mcm5l1f_cf_w_0_170_s_0_225=4.94e-12
.param mcm5l1f_ca_w_0_170_s_0_270=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_270=5.92e-11
.param mcm5l1f_cf_w_0_170_s_0_270=5.86e-12
.param mcm5l1f_ca_w_0_170_s_0_360=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_360=4.80e-11
.param mcm5l1f_cf_w_0_170_s_0_360=7.86e-12
.param mcm5l1f_ca_w_0_170_s_0_450=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_450=4.09e-11
.param mcm5l1f_cf_w_0_170_s_0_450=9.44e-12
.param mcm5l1f_ca_w_0_170_s_0_540=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_540=3.52e-11
.param mcm5l1f_cf_w_0_170_s_0_540=1.13e-11
.param mcm5l1f_ca_w_0_170_s_0_720=4.49e-05
.param mcm5l1f_cc_w_0_170_s_0_720=2.77e-11
.param mcm5l1f_cf_w_0_170_s_0_720=1.43e-11
.param mcm5l1f_ca_w_0_170_s_1_080=4.49e-05
.param mcm5l1f_cc_w_0_170_s_1_080=1.85e-11
.param mcm5l1f_cf_w_0_170_s_1_080=1.94e-11
.param mcm5l1f_ca_w_0_170_s_1_980=4.49e-05
.param mcm5l1f_cc_w_0_170_s_1_980=8.13e-12
.param mcm5l1f_cf_w_0_170_s_1_980=2.70e-11
.param mcm5l1f_ca_w_0_170_s_4_500=4.49e-05
.param mcm5l1f_cc_w_0_170_s_4_500=1.29e-12
.param mcm5l1f_cf_w_0_170_s_4_500=3.31e-11
.param mcm5l1f_ca_w_1_360_s_0_180=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_180=9.67e-11
.param mcm5l1f_cf_w_1_360_s_0_180=3.97e-12
.param mcm5l1f_ca_w_1_360_s_0_225=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_225=8.35e-11
.param mcm5l1f_cf_w_1_360_s_0_225=4.93e-12
.param mcm5l1f_ca_w_1_360_s_0_270=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_270=7.42e-11
.param mcm5l1f_cf_w_1_360_s_0_270=5.87e-12
.param mcm5l1f_ca_w_1_360_s_0_360=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_360=6.12e-11
.param mcm5l1f_cf_w_1_360_s_0_360=7.72e-12
.param mcm5l1f_ca_w_1_360_s_0_450=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_450=5.24e-11
.param mcm5l1f_cf_w_1_360_s_0_450=9.51e-12
.param mcm5l1f_ca_w_1_360_s_0_540=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_540=4.59e-11
.param mcm5l1f_cf_w_1_360_s_0_540=1.12e-11
.param mcm5l1f_ca_w_1_360_s_0_720=4.49e-05
.param mcm5l1f_cc_w_1_360_s_0_720=3.67e-11
.param mcm5l1f_cf_w_1_360_s_0_720=1.44e-11
.param mcm5l1f_ca_w_1_360_s_1_080=4.49e-05
.param mcm5l1f_cc_w_1_360_s_1_080=2.53e-11
.param mcm5l1f_cf_w_1_360_s_1_080=1.98e-11
.param mcm5l1f_ca_w_1_360_s_1_980=4.49e-05
.param mcm5l1f_cc_w_1_360_s_1_980=1.20e-11
.param mcm5l1f_cf_w_1_360_s_1_980=2.90e-11
.param mcm5l1f_ca_w_1_360_s_4_500=4.49e-05
.param mcm5l1f_cc_w_1_360_s_4_500=2.14e-12
.param mcm5l1f_cf_w_1_360_s_4_500=3.76e-11
.param mcm5l1d_ca_w_0_170_s_0_180=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_180=7.65e-11
.param mcm5l1d_cf_w_0_170_s_0_180=5.54e-12
.param mcm5l1d_ca_w_0_170_s_0_225=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_225=6.45e-11
.param mcm5l1d_cf_w_0_170_s_0_225=6.86e-12
.param mcm5l1d_ca_w_0_170_s_0_270=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_270=5.64e-11
.param mcm5l1d_cf_w_0_170_s_0_270=8.13e-12
.param mcm5l1d_ca_w_0_170_s_0_360=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_360=4.49e-11
.param mcm5l1d_cf_w_0_170_s_0_360=1.08e-11
.param mcm5l1d_ca_w_0_170_s_0_450=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_450=3.77e-11
.param mcm5l1d_cf_w_0_170_s_0_450=1.29e-11
.param mcm5l1d_ca_w_0_170_s_0_540=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_540=3.18e-11
.param mcm5l1d_cf_w_0_170_s_0_540=1.53e-11
.param mcm5l1d_ca_w_0_170_s_0_720=6.33e-05
.param mcm5l1d_cc_w_0_170_s_0_720=2.41e-11
.param mcm5l1d_cf_w_0_170_s_0_720=1.91e-11
.param mcm5l1d_ca_w_0_170_s_1_080=6.33e-05
.param mcm5l1d_cc_w_0_170_s_1_080=1.51e-11
.param mcm5l1d_cf_w_0_170_s_1_080=2.50e-11
.param mcm5l1d_ca_w_0_170_s_1_980=6.33e-05
.param mcm5l1d_cc_w_0_170_s_1_980=5.84e-12
.param mcm5l1d_cf_w_0_170_s_1_980=3.25e-11
.param mcm5l1d_ca_w_0_170_s_4_500=6.33e-05
.param mcm5l1d_cc_w_0_170_s_4_500=7.85e-13
.param mcm5l1d_cf_w_0_170_s_4_500=3.72e-11
.param mcm5l1d_ca_w_1_360_s_0_180=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_180=9.23e-11
.param mcm5l1d_cf_w_1_360_s_0_180=5.53e-12
.param mcm5l1d_ca_w_1_360_s_0_225=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_225=7.91e-11
.param mcm5l1d_cf_w_1_360_s_0_225=6.86e-12
.param mcm5l1d_ca_w_1_360_s_0_270=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_270=6.98e-11
.param mcm5l1d_cf_w_1_360_s_0_270=8.15e-12
.param mcm5l1d_ca_w_1_360_s_0_360=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_360=5.68e-11
.param mcm5l1d_cf_w_1_360_s_0_360=1.06e-11
.param mcm5l1d_ca_w_1_360_s_0_450=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_450=4.81e-11
.param mcm5l1d_cf_w_1_360_s_0_450=1.30e-11
.param mcm5l1d_ca_w_1_360_s_0_540=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_540=4.16e-11
.param mcm5l1d_cf_w_1_360_s_0_540=1.52e-11
.param mcm5l1d_ca_w_1_360_s_0_720=6.33e-05
.param mcm5l1d_cc_w_1_360_s_0_720=3.25e-11
.param mcm5l1d_cf_w_1_360_s_0_720=1.92e-11
.param mcm5l1d_ca_w_1_360_s_1_080=6.33e-05
.param mcm5l1d_cc_w_1_360_s_1_080=2.14e-11
.param mcm5l1d_cf_w_1_360_s_1_080=2.56e-11
.param mcm5l1d_ca_w_1_360_s_1_980=6.33e-05
.param mcm5l1d_cc_w_1_360_s_1_980=9.30e-12
.param mcm5l1d_cf_w_1_360_s_1_980=3.51e-11
.param mcm5l1d_ca_w_1_360_s_4_500=6.33e-05
.param mcm5l1d_cc_w_1_360_s_4_500=1.49e-12
.param mcm5l1d_cf_w_1_360_s_4_500=4.23e-11
.param mcm5l1p1_ca_w_0_170_s_0_180=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_180=7.21e-11
.param mcm5l1p1_cf_w_0_170_s_0_180=8.78e-12
.param mcm5l1p1_ca_w_0_170_s_0_225=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_225=6.01e-11
.param mcm5l1p1_cf_w_0_170_s_0_225=1.08e-11
.param mcm5l1p1_ca_w_0_170_s_0_270=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_270=5.17e-11
.param mcm5l1p1_cf_w_0_170_s_0_270=1.27e-11
.param mcm5l1p1_ca_w_0_170_s_0_360=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_360=4.00e-11
.param mcm5l1p1_cf_w_0_170_s_0_360=1.66e-11
.param mcm5l1p1_ca_w_0_170_s_0_450=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_450=3.27e-11
.param mcm5l1p1_cf_w_0_170_s_0_450=1.96e-11
.param mcm5l1p1_ca_w_0_170_s_0_540=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_540=2.68e-11
.param mcm5l1p1_cf_w_0_170_s_0_540=2.28e-11
.param mcm5l1p1_ca_w_0_170_s_0_720=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_0_720=1.92e-11
.param mcm5l1p1_cf_w_0_170_s_0_720=2.76e-11
.param mcm5l1p1_ca_w_0_170_s_1_080=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_1_080=1.09e-11
.param mcm5l1p1_cf_w_0_170_s_1_080=3.40e-11
.param mcm5l1p1_ca_w_0_170_s_1_980=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_1_980=3.61e-12
.param mcm5l1p1_cf_w_0_170_s_1_980=4.05e-11
.param mcm5l1p1_ca_w_0_170_s_4_500=1.02e-04
.param mcm5l1p1_cc_w_0_170_s_4_500=4.47e-13
.param mcm5l1p1_cf_w_0_170_s_4_500=4.35e-11
.param mcm5l1p1_ca_w_1_360_s_0_180=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_180=8.63e-11
.param mcm5l1p1_cf_w_1_360_s_0_180=8.86e-12
.param mcm5l1p1_ca_w_1_360_s_0_225=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_225=7.34e-11
.param mcm5l1p1_cf_w_1_360_s_0_225=1.09e-11
.param mcm5l1p1_ca_w_1_360_s_0_270=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_270=6.39e-11
.param mcm5l1p1_cf_w_1_360_s_0_270=1.28e-11
.param mcm5l1p1_ca_w_1_360_s_0_360=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_360=5.11e-11
.param mcm5l1p1_cf_w_1_360_s_0_360=1.65e-11
.param mcm5l1p1_ca_w_1_360_s_0_450=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_450=4.24e-11
.param mcm5l1p1_cf_w_1_360_s_0_450=1.98e-11
.param mcm5l1p1_ca_w_1_360_s_0_540=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_540=3.60e-11
.param mcm5l1p1_cf_w_1_360_s_0_540=2.28e-11
.param mcm5l1p1_ca_w_1_360_s_0_720=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_0_720=2.72e-11
.param mcm5l1p1_cf_w_1_360_s_0_720=2.79e-11
.param mcm5l1p1_ca_w_1_360_s_1_080=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_1_080=1.70e-11
.param mcm5l1p1_cf_w_1_360_s_1_080=3.53e-11
.param mcm5l1p1_ca_w_1_360_s_1_980=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_1_980=6.69e-12
.param mcm5l1p1_cf_w_1_360_s_1_980=4.41e-11
.param mcm5l1p1_ca_w_1_360_s_4_500=1.02e-04
.param mcm5l1p1_cc_w_1_360_s_4_500=9.85e-13
.param mcm5l1p1_cf_w_1_360_s_4_500=4.96e-11
.param mcrdll1f_ca_w_0_170_s_0_180=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_180=7.95e-11
.param mcrdll1f_cf_w_0_170_s_0_180=3.51e-12
.param mcrdll1f_ca_w_0_170_s_0_225=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_225=6.78e-11
.param mcrdll1f_cf_w_0_170_s_0_225=4.35e-12
.param mcrdll1f_ca_w_0_170_s_0_270=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_270=6.01e-11
.param mcrdll1f_cf_w_0_170_s_0_270=5.18e-12
.param mcrdll1f_ca_w_0_170_s_0_360=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_360=4.91e-11
.param mcrdll1f_cf_w_0_170_s_0_360=6.97e-12
.param mcrdll1f_ca_w_0_170_s_0_450=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_450=4.22e-11
.param mcrdll1f_cf_w_0_170_s_0_450=8.36e-12
.param mcrdll1f_ca_w_0_170_s_0_540=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_540=3.66e-11
.param mcrdll1f_cf_w_0_170_s_0_540=1.01e-11
.param mcrdll1f_ca_w_0_170_s_0_720=3.97e-05
.param mcrdll1f_cc_w_0_170_s_0_720=2.92e-11
.param mcrdll1f_cf_w_0_170_s_0_720=1.28e-11
.param mcrdll1f_ca_w_0_170_s_1_080=3.97e-05
.param mcrdll1f_cc_w_0_170_s_1_080=2.03e-11
.param mcrdll1f_cf_w_0_170_s_1_080=1.76e-11
.param mcrdll1f_ca_w_0_170_s_1_980=3.97e-05
.param mcrdll1f_cc_w_0_170_s_1_980=1.02e-11
.param mcrdll1f_cf_w_0_170_s_1_980=2.49e-11
.param mcrdll1f_ca_w_0_170_s_4_500=3.97e-05
.param mcrdll1f_cc_w_0_170_s_4_500=2.50e-12
.param mcrdll1f_cf_w_0_170_s_4_500=3.18e-11
.param mcrdll1f_ca_w_1_360_s_0_180=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_180=1.00e-10
.param mcrdll1f_cf_w_1_360_s_0_180=3.51e-12
.param mcrdll1f_ca_w_1_360_s_0_225=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_225=8.69e-11
.param mcrdll1f_cf_w_1_360_s_0_225=4.36e-12
.param mcrdll1f_ca_w_1_360_s_0_270=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_270=7.76e-11
.param mcrdll1f_cf_w_1_360_s_0_270=5.19e-12
.param mcrdll1f_ca_w_1_360_s_0_360=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_360=6.49e-11
.param mcrdll1f_cf_w_1_360_s_0_360=6.83e-12
.param mcrdll1f_ca_w_1_360_s_0_450=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_450=5.63e-11
.param mcrdll1f_cf_w_1_360_s_0_450=8.42e-12
.param mcrdll1f_ca_w_1_360_s_0_540=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_540=4.98e-11
.param mcrdll1f_cf_w_1_360_s_0_540=9.94e-12
.param mcrdll1f_ca_w_1_360_s_0_720=3.97e-05
.param mcrdll1f_cc_w_1_360_s_0_720=4.08e-11
.param mcrdll1f_cf_w_1_360_s_0_720=1.28e-11
.param mcrdll1f_ca_w_1_360_s_1_080=3.97e-05
.param mcrdll1f_cc_w_1_360_s_1_080=2.98e-11
.param mcrdll1f_cf_w_1_360_s_1_080=1.78e-11
.param mcrdll1f_ca_w_1_360_s_1_980=3.97e-05
.param mcrdll1f_cc_w_1_360_s_1_980=1.63e-11
.param mcrdll1f_cf_w_1_360_s_1_980=2.67e-11
.param mcrdll1f_ca_w_1_360_s_4_500=3.97e-05
.param mcrdll1f_cc_w_1_360_s_4_500=4.82e-12
.param mcrdll1f_cf_w_1_360_s_4_500=3.66e-11
.param mcrdll1d_ca_w_0_170_s_0_180=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_180=7.71e-11
.param mcrdll1d_cf_w_0_170_s_0_180=5.08e-12
.param mcrdll1d_ca_w_0_170_s_0_225=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_225=6.53e-11
.param mcrdll1d_cf_w_0_170_s_0_225=6.29e-12
.param mcrdll1d_ca_w_0_170_s_0_270=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_270=5.73e-11
.param mcrdll1d_cf_w_0_170_s_0_270=7.44e-12
.param mcrdll1d_ca_w_0_170_s_0_360=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_360=4.60e-11
.param mcrdll1d_cf_w_0_170_s_0_360=9.92e-12
.param mcrdll1d_ca_w_0_170_s_0_450=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_450=3.89e-11
.param mcrdll1d_cf_w_0_170_s_0_450=1.19e-11
.param mcrdll1d_ca_w_0_170_s_0_540=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_540=3.32e-11
.param mcrdll1d_cf_w_0_170_s_0_540=1.41e-11
.param mcrdll1d_ca_w_0_170_s_0_720=5.80e-05
.param mcrdll1d_cc_w_0_170_s_0_720=2.56e-11
.param mcrdll1d_cf_w_0_170_s_0_720=1.77e-11
.param mcrdll1d_ca_w_0_170_s_1_080=5.80e-05
.param mcrdll1d_cc_w_0_170_s_1_080=1.67e-11
.param mcrdll1d_cf_w_0_170_s_1_080=2.34e-11
.param mcrdll1d_ca_w_0_170_s_1_980=5.80e-05
.param mcrdll1d_cc_w_0_170_s_1_980=7.48e-12
.param mcrdll1d_cf_w_0_170_s_1_980=3.09e-11
.param mcrdll1d_ca_w_0_170_s_4_500=5.80e-05
.param mcrdll1d_cc_w_0_170_s_4_500=1.61e-12
.param mcrdll1d_cf_w_0_170_s_4_500=3.64e-11
.param mcrdll1d_ca_w_1_360_s_0_180=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_180=9.55e-11
.param mcrdll1d_cf_w_1_360_s_0_180=5.08e-12
.param mcrdll1d_ca_w_1_360_s_0_225=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_225=8.26e-11
.param mcrdll1d_cf_w_1_360_s_0_225=6.29e-12
.param mcrdll1d_ca_w_1_360_s_0_270=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_270=7.32e-11
.param mcrdll1d_cf_w_1_360_s_0_270=7.47e-12
.param mcrdll1d_ca_w_1_360_s_0_360=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_360=6.05e-11
.param mcrdll1d_cf_w_1_360_s_0_360=9.77e-12
.param mcrdll1d_ca_w_1_360_s_0_450=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_450=5.19e-11
.param mcrdll1d_cf_w_1_360_s_0_450=1.19e-11
.param mcrdll1d_ca_w_1_360_s_0_540=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_540=4.55e-11
.param mcrdll1d_cf_w_1_360_s_0_540=1.40e-11
.param mcrdll1d_ca_w_1_360_s_0_720=5.80e-05
.param mcrdll1d_cc_w_1_360_s_0_720=3.65e-11
.param mcrdll1d_cf_w_1_360_s_0_720=1.78e-11
.param mcrdll1d_ca_w_1_360_s_1_080=5.80e-05
.param mcrdll1d_cc_w_1_360_s_1_080=2.56e-11
.param mcrdll1d_cf_w_1_360_s_1_080=2.39e-11
.param mcrdll1d_ca_w_1_360_s_1_980=5.80e-05
.param mcrdll1d_cc_w_1_360_s_1_980=1.31e-11
.param mcrdll1d_cf_w_1_360_s_1_980=3.34e-11
.param mcrdll1d_ca_w_1_360_s_4_500=5.80e-05
.param mcrdll1d_cc_w_1_360_s_4_500=3.58e-12
.param mcrdll1d_cf_w_1_360_s_4_500=4.22e-11
.param mcrdll1p1_ca_w_0_170_s_0_180=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_180=7.29e-11
.param mcrdll1p1_cf_w_0_170_s_0_180=8.32e-12
.param mcrdll1p1_ca_w_0_170_s_0_225=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_225=6.09e-11
.param mcrdll1p1_cf_w_0_170_s_0_225=1.02e-11
.param mcrdll1p1_ca_w_0_170_s_0_270=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_270=5.27e-11
.param mcrdll1p1_cf_w_0_170_s_0_270=1.20e-11
.param mcrdll1p1_ca_w_0_170_s_0_360=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_360=4.10e-11
.param mcrdll1p1_cf_w_0_170_s_0_360=1.58e-11
.param mcrdll1p1_ca_w_0_170_s_0_450=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_450=3.39e-11
.param mcrdll1p1_cf_w_0_170_s_0_450=1.86e-11
.param mcrdll1p1_ca_w_0_170_s_0_540=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_540=2.80e-11
.param mcrdll1p1_cf_w_0_170_s_0_540=2.17e-11
.param mcrdll1p1_ca_w_0_170_s_0_720=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_0_720=2.05e-11
.param mcrdll1p1_cf_w_0_170_s_0_720=2.64e-11
.param mcrdll1p1_ca_w_0_170_s_1_080=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_1_080=1.21e-11
.param mcrdll1p1_cf_w_0_170_s_1_080=3.28e-11
.param mcrdll1p1_ca_w_0_170_s_1_980=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_1_980=4.79e-12
.param mcrdll1p1_cf_w_0_170_s_1_980=3.95e-11
.param mcrdll1p1_ca_w_0_170_s_4_500=9.69e-05
.param mcrdll1p1_cc_w_0_170_s_4_500=9.61e-13
.param mcrdll1p1_cf_w_0_170_s_4_500=4.32e-11
.param mcrdll1p1_ca_w_1_360_s_0_180=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_180=8.97e-11
.param mcrdll1p1_cf_w_1_360_s_0_180=8.41e-12
.param mcrdll1p1_ca_w_1_360_s_0_225=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_225=7.67e-11
.param mcrdll1p1_cf_w_1_360_s_0_225=1.03e-11
.param mcrdll1p1_ca_w_1_360_s_0_270=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_270=6.74e-11
.param mcrdll1p1_cf_w_1_360_s_0_270=1.22e-11
.param mcrdll1p1_ca_w_1_360_s_0_360=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_360=5.46e-11
.param mcrdll1p1_cf_w_1_360_s_0_360=1.56e-11
.param mcrdll1p1_ca_w_1_360_s_0_450=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_450=4.61e-11
.param mcrdll1p1_cf_w_1_360_s_0_450=1.88e-11
.param mcrdll1p1_ca_w_1_360_s_0_540=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_540=3.98e-11
.param mcrdll1p1_cf_w_1_360_s_0_540=2.17e-11
.param mcrdll1p1_ca_w_1_360_s_0_720=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_0_720=3.11e-11
.param mcrdll1p1_cf_w_1_360_s_0_720=2.67e-11
.param mcrdll1p1_ca_w_1_360_s_1_080=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_1_080=2.09e-11
.param mcrdll1p1_cf_w_1_360_s_1_080=3.39e-11
.param mcrdll1p1_ca_w_1_360_s_1_980=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_1_980=9.91e-12
.param mcrdll1p1_cf_w_1_360_s_1_980=4.34e-11
.param mcrdll1p1_ca_w_1_360_s_4_500=9.69e-05
.param mcrdll1p1_cc_w_1_360_s_4_500=2.56e-12
.param mcrdll1p1_cf_w_1_360_s_4_500=5.04e-11
.param mcm2m1f_ca_w_0_140_s_0_140=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_140=9.21e-11
.param mcm2m1f_cf_w_0_140_s_0_140=9.79e-12
.param mcm2m1f_ca_w_0_140_s_0_175=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_175=9.00e-11
.param mcm2m1f_cf_w_0_140_s_0_175=1.20e-11
.param mcm2m1f_ca_w_0_140_s_0_210=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_210=8.45e-11
.param mcm2m1f_cf_w_0_140_s_0_210=1.42e-11
.param mcm2m1f_ca_w_0_140_s_0_280=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_280=7.12e-11
.param mcm2m1f_cf_w_0_140_s_0_280=1.84e-11
.param mcm2m1f_ca_w_0_140_s_0_350=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_350=5.93e-11
.param mcm2m1f_cf_w_0_140_s_0_350=2.23e-11
.param mcm2m1f_ca_w_0_140_s_0_420=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_420=4.91e-11
.param mcm2m1f_cf_w_0_140_s_0_420=2.61e-11
.param mcm2m1f_ca_w_0_140_s_0_560=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_560=3.50e-11
.param mcm2m1f_cf_w_0_140_s_0_560=3.22e-11
.param mcm2m1f_ca_w_0_140_s_0_840=1.54e-04
.param mcm2m1f_cc_w_0_140_s_0_840=1.97e-11
.param mcm2m1f_cf_w_0_140_s_0_840=4.17e-11
.param mcm2m1f_ca_w_0_140_s_1_540=1.54e-04
.param mcm2m1f_cc_w_0_140_s_1_540=5.79e-12
.param mcm2m1f_cf_w_0_140_s_1_540=5.32e-11
.param mcm2m1f_ca_w_0_140_s_3_500=1.54e-04
.param mcm2m1f_cc_w_0_140_s_3_500=3.20e-13
.param mcm2m1f_cf_w_0_140_s_3_500=5.86e-11
.param mcm2m1f_ca_w_1_120_s_0_140=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_140=1.01e-10
.param mcm2m1f_cf_w_1_120_s_0_140=9.82e-12
.param mcm2m1f_ca_w_1_120_s_0_175=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_175=9.83e-11
.param mcm2m1f_cf_w_1_120_s_0_175=1.21e-11
.param mcm2m1f_ca_w_1_120_s_0_210=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_210=9.13e-11
.param mcm2m1f_cf_w_1_120_s_0_210=1.43e-11
.param mcm2m1f_ca_w_1_120_s_0_280=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_280=7.75e-11
.param mcm2m1f_cf_w_1_120_s_0_280=1.84e-11
.param mcm2m1f_ca_w_1_120_s_0_350=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_350=6.48e-11
.param mcm2m1f_cf_w_1_120_s_0_350=2.24e-11
.param mcm2m1f_ca_w_1_120_s_0_420=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_420=5.39e-11
.param mcm2m1f_cf_w_1_120_s_0_420=2.61e-11
.param mcm2m1f_ca_w_1_120_s_0_560=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_560=3.86e-11
.param mcm2m1f_cf_w_1_120_s_0_560=3.25e-11
.param mcm2m1f_ca_w_1_120_s_0_840=1.54e-04
.param mcm2m1f_cc_w_1_120_s_0_840=2.21e-11
.param mcm2m1f_cf_w_1_120_s_0_840=4.21e-11
.param mcm2m1f_ca_w_1_120_s_1_540=1.54e-04
.param mcm2m1f_cc_w_1_120_s_1_540=6.77e-12
.param mcm2m1f_cf_w_1_120_s_1_540=5.43e-11
.param mcm2m1f_ca_w_1_120_s_3_500=1.54e-04
.param mcm2m1f_cc_w_1_120_s_3_500=3.65e-13
.param mcm2m1f_cf_w_1_120_s_3_500=6.08e-11
.param mcm2m1d_ca_w_0_140_s_0_140=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_140=9.13e-11
.param mcm2m1d_cf_w_0_140_s_0_140=1.03e-11
.param mcm2m1d_ca_w_0_140_s_0_175=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_175=8.90e-11
.param mcm2m1d_cf_w_0_140_s_0_175=1.27e-11
.param mcm2m1d_ca_w_0_140_s_0_210=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_210=8.32e-11
.param mcm2m1d_cf_w_0_140_s_0_210=1.50e-11
.param mcm2m1d_ca_w_0_140_s_0_280=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_280=6.98e-11
.param mcm2m1d_cf_w_0_140_s_0_280=1.95e-11
.param mcm2m1d_ca_w_0_140_s_0_350=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_350=5.79e-11
.param mcm2m1d_cf_w_0_140_s_0_350=2.36e-11
.param mcm2m1d_ca_w_0_140_s_0_420=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_420=4.76e-11
.param mcm2m1d_cf_w_0_140_s_0_420=2.76e-11
.param mcm2m1d_ca_w_0_140_s_0_560=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_560=3.33e-11
.param mcm2m1d_cf_w_0_140_s_0_560=3.41e-11
.param mcm2m1d_ca_w_0_140_s_0_840=1.62e-04
.param mcm2m1d_cc_w_0_140_s_0_840=1.78e-11
.param mcm2m1d_cf_w_0_140_s_0_840=4.39e-11
.param mcm2m1d_ca_w_0_140_s_1_540=1.62e-04
.param mcm2m1d_cc_w_0_140_s_1_540=4.57e-12
.param mcm2m1d_cf_w_0_140_s_1_540=5.53e-11
.param mcm2m1d_ca_w_0_140_s_3_500=1.62e-04
.param mcm2m1d_cc_w_0_140_s_3_500=1.75e-13
.param mcm2m1d_cf_w_0_140_s_3_500=5.99e-11
.param mcm2m1d_ca_w_1_120_s_0_140=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_140=9.89e-11
.param mcm2m1d_cf_w_1_120_s_0_140=1.04e-11
.param mcm2m1d_ca_w_1_120_s_0_175=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_175=9.56e-11
.param mcm2m1d_cf_w_1_120_s_0_175=1.28e-11
.param mcm2m1d_ca_w_1_120_s_0_210=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_210=8.86e-11
.param mcm2m1d_cf_w_1_120_s_0_210=1.51e-11
.param mcm2m1d_ca_w_1_120_s_0_280=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_280=7.49e-11
.param mcm2m1d_cf_w_1_120_s_0_280=1.95e-11
.param mcm2m1d_ca_w_1_120_s_0_350=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_350=6.19e-11
.param mcm2m1d_cf_w_1_120_s_0_350=2.37e-11
.param mcm2m1d_ca_w_1_120_s_0_420=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_420=5.10e-11
.param mcm2m1d_cf_w_1_120_s_0_420=2.76e-11
.param mcm2m1d_ca_w_1_120_s_0_560=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_560=3.58e-11
.param mcm2m1d_cf_w_1_120_s_0_560=3.44e-11
.param mcm2m1d_ca_w_1_120_s_0_840=1.62e-04
.param mcm2m1d_cc_w_1_120_s_0_840=1.95e-11
.param mcm2m1d_cf_w_1_120_s_0_840=4.44e-11
.param mcm2m1d_ca_w_1_120_s_1_540=1.62e-04
.param mcm2m1d_cc_w_1_120_s_1_540=5.09e-12
.param mcm2m1d_cf_w_1_120_s_1_540=5.64e-11
.param mcm2m1d_ca_w_1_120_s_3_500=1.62e-04
.param mcm2m1d_cc_w_1_120_s_3_500=1.70e-13
.param mcm2m1d_cf_w_1_120_s_3_500=6.15e-11
.param mcm2m1p1_ca_w_0_140_s_0_140=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_140=9.03e-11
.param mcm2m1p1_cf_w_0_140_s_0_140=1.11e-11
.param mcm2m1p1_ca_w_0_140_s_0_175=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_175=8.77e-11
.param mcm2m1p1_cf_w_0_140_s_0_175=1.37e-11
.param mcm2m1p1_ca_w_0_140_s_0_210=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_210=8.13e-11
.param mcm2m1p1_cf_w_0_140_s_0_210=1.62e-11
.param mcm2m1p1_ca_w_0_140_s_0_280=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_280=6.80e-11
.param mcm2m1p1_cf_w_0_140_s_0_280=2.10e-11
.param mcm2m1p1_ca_w_0_140_s_0_350=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_350=5.59e-11
.param mcm2m1p1_cf_w_0_140_s_0_350=2.54e-11
.param mcm2m1p1_ca_w_0_140_s_0_420=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_420=4.55e-11
.param mcm2m1p1_cf_w_0_140_s_0_420=2.97e-11
.param mcm2m1p1_ca_w_0_140_s_0_560=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_560=3.09e-11
.param mcm2m1p1_cf_w_0_140_s_0_560=3.67e-11
.param mcm2m1p1_ca_w_0_140_s_0_840=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_0_840=1.56e-11
.param mcm2m1p1_cf_w_0_140_s_0_840=4.70e-11
.param mcm2m1p1_ca_w_0_140_s_1_540=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_1_540=3.31e-12
.param mcm2m1p1_cf_w_0_140_s_1_540=5.80e-11
.param mcm2m1p1_ca_w_0_140_s_3_500=1.73e-04
.param mcm2m1p1_cc_w_0_140_s_3_500=1.25e-13
.param mcm2m1p1_cf_w_0_140_s_3_500=6.16e-11
.param mcm2m1p1_ca_w_1_120_s_0_140=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_140=9.55e-11
.param mcm2m1p1_cf_w_1_120_s_0_140=1.12e-11
.param mcm2m1p1_ca_w_1_120_s_0_175=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_175=9.24e-11
.param mcm2m1p1_cf_w_1_120_s_0_175=1.38e-11
.param mcm2m1p1_ca_w_1_120_s_0_210=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_210=8.64e-11
.param mcm2m1p1_cf_w_1_120_s_0_210=1.63e-11
.param mcm2m1p1_ca_w_1_120_s_0_280=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_280=7.16e-11
.param mcm2m1p1_cf_w_1_120_s_0_280=2.11e-11
.param mcm2m1p1_ca_w_1_120_s_0_350=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_350=5.87e-11
.param mcm2m1p1_cf_w_1_120_s_0_350=2.56e-11
.param mcm2m1p1_ca_w_1_120_s_0_420=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_420=4.79e-11
.param mcm2m1p1_cf_w_1_120_s_0_420=2.98e-11
.param mcm2m1p1_ca_w_1_120_s_0_560=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_560=3.25e-11
.param mcm2m1p1_cf_w_1_120_s_0_560=3.70e-11
.param mcm2m1p1_ca_w_1_120_s_0_840=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_0_840=1.66e-11
.param mcm2m1p1_cf_w_1_120_s_0_840=4.75e-11
.param mcm2m1p1_ca_w_1_120_s_1_540=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_1_540=3.54e-12
.param mcm2m1p1_cf_w_1_120_s_1_540=5.88e-11
.param mcm2m1p1_ca_w_1_120_s_3_500=1.73e-04
.param mcm2m1p1_cc_w_1_120_s_3_500=1.20e-13
.param mcm2m1p1_cf_w_1_120_s_3_500=6.28e-11
.param mcm2m1l1_ca_w_0_140_s_0_140=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_140=8.35e-11
.param mcm2m1l1_cf_w_0_140_s_0_140=1.54e-11
.param mcm2m1l1_ca_w_0_140_s_0_175=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_175=8.06e-11
.param mcm2m1l1_cf_w_0_140_s_0_175=1.92e-11
.param mcm2m1l1_ca_w_0_140_s_0_210=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_210=7.38e-11
.param mcm2m1l1_cf_w_0_140_s_0_210=2.28e-11
.param mcm2m1l1_ca_w_0_140_s_0_280=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_280=6.02e-11
.param mcm2m1l1_cf_w_0_140_s_0_280=2.96e-11
.param mcm2m1l1_ca_w_0_140_s_0_350=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_350=4.74e-11
.param mcm2m1l1_cf_w_0_140_s_0_350=3.60e-11
.param mcm2m1l1_ca_w_0_140_s_0_420=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_420=3.68e-11
.param mcm2m1l1_cf_w_0_140_s_0_420=4.16e-11
.param mcm2m1l1_ca_w_0_140_s_0_560=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_560=2.26e-11
.param mcm2m1l1_cf_w_0_140_s_0_560=5.08e-11
.param mcm2m1l1_ca_w_0_140_s_0_840=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_0_840=8.81e-12
.param mcm2m1l1_cf_w_0_140_s_0_840=6.23e-11
.param mcm2m1l1_ca_w_0_140_s_1_540=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_1_540=9.45e-13
.param mcm2m1l1_cf_w_0_140_s_1_540=7.06e-11
.param mcm2m1l1_ca_w_0_140_s_3_500=2.42e-04
.param mcm2m1l1_cc_w_0_140_s_3_500=2.50e-14
.param mcm2m1l1_cf_w_0_140_s_3_500=7.20e-11
.param mcm2m1l1_ca_w_1_120_s_0_140=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_140=8.49e-11
.param mcm2m1l1_cf_w_1_120_s_0_140=1.55e-11
.param mcm2m1l1_ca_w_1_120_s_0_175=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_175=8.16e-11
.param mcm2m1l1_cf_w_1_120_s_0_175=1.93e-11
.param mcm2m1l1_ca_w_1_120_s_0_210=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_210=7.54e-11
.param mcm2m1l1_cf_w_1_120_s_0_210=2.29e-11
.param mcm2m1l1_ca_w_1_120_s_0_280=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_280=6.07e-11
.param mcm2m1l1_cf_w_1_120_s_0_280=2.97e-11
.param mcm2m1l1_ca_w_1_120_s_0_350=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_350=4.79e-11
.param mcm2m1l1_cf_w_1_120_s_0_350=3.60e-11
.param mcm2m1l1_ca_w_1_120_s_0_420=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_420=3.72e-11
.param mcm2m1l1_cf_w_1_120_s_0_420=4.17e-11
.param mcm2m1l1_ca_w_1_120_s_0_560=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_560=2.28e-11
.param mcm2m1l1_cf_w_1_120_s_0_560=5.10e-11
.param mcm2m1l1_ca_w_1_120_s_0_840=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_0_840=9.00e-12
.param mcm2m1l1_cf_w_1_120_s_0_840=6.26e-11
.param mcm2m1l1_ca_w_1_120_s_1_540=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_1_540=9.50e-13
.param mcm2m1l1_cf_w_1_120_s_1_540=7.09e-11
.param mcm2m1l1_ca_w_1_120_s_3_500=2.42e-04
.param mcm2m1l1_cc_w_1_120_s_3_500=5.00e-14
.param mcm2m1l1_cf_w_1_120_s_3_500=7.24e-11
.param mcm3m1f_ca_w_0_140_s_0_140=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_140=1.01e-10
.param mcm3m1f_cf_w_0_140_s_0_140=4.03e-12
.param mcm3m1f_ca_w_0_140_s_0_175=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_175=9.91e-11
.param mcm3m1f_cf_w_0_140_s_0_175=5.02e-12
.param mcm3m1f_ca_w_0_140_s_0_210=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_210=9.37e-11
.param mcm3m1f_cf_w_0_140_s_0_210=6.02e-12
.param mcm3m1f_ca_w_0_140_s_0_280=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_280=8.17e-11
.param mcm3m1f_cf_w_0_140_s_0_280=7.95e-12
.param mcm3m1f_ca_w_0_140_s_0_350=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_350=7.03e-11
.param mcm3m1f_cf_w_0_140_s_0_350=9.85e-12
.param mcm3m1f_ca_w_0_140_s_0_420=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_420=5.99e-11
.param mcm3m1f_cf_w_0_140_s_0_420=1.18e-11
.param mcm3m1f_ca_w_0_140_s_0_560=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_560=4.61e-11
.param mcm3m1f_cf_w_0_140_s_0_560=1.52e-11
.param mcm3m1f_ca_w_0_140_s_0_840=5.87e-05
.param mcm3m1f_cc_w_0_140_s_0_840=3.00e-11
.param mcm3m1f_cf_w_0_140_s_0_840=2.14e-11
.param mcm3m1f_ca_w_0_140_s_1_540=5.87e-05
.param mcm3m1f_cc_w_0_140_s_1_540=1.25e-11
.param mcm3m1f_cf_w_0_140_s_1_540=3.23e-11
.param mcm3m1f_ca_w_0_140_s_3_500=5.87e-05
.param mcm3m1f_cc_w_0_140_s_3_500=1.40e-12
.param mcm3m1f_cf_w_0_140_s_3_500=4.19e-11
.param mcm3m1f_ca_w_1_120_s_0_140=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_140=1.16e-10
.param mcm3m1f_cf_w_1_120_s_0_140=4.06e-12
.param mcm3m1f_ca_w_1_120_s_0_175=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_175=1.13e-10
.param mcm3m1f_cf_w_1_120_s_0_175=5.06e-12
.param mcm3m1f_ca_w_1_120_s_0_210=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_210=1.06e-10
.param mcm3m1f_cf_w_1_120_s_0_210=6.05e-12
.param mcm3m1f_ca_w_1_120_s_0_280=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_280=9.17e-11
.param mcm3m1f_cf_w_1_120_s_0_280=7.99e-12
.param mcm3m1f_ca_w_1_120_s_0_350=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_350=7.90e-11
.param mcm3m1f_cf_w_1_120_s_0_350=9.92e-12
.param mcm3m1f_ca_w_1_120_s_0_420=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_420=6.80e-11
.param mcm3m1f_cf_w_1_120_s_0_420=1.18e-11
.param mcm3m1f_ca_w_1_120_s_0_560=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_560=5.21e-11
.param mcm3m1f_cf_w_1_120_s_0_560=1.54e-11
.param mcm3m1f_ca_w_1_120_s_0_840=5.87e-05
.param mcm3m1f_cc_w_1_120_s_0_840=3.39e-11
.param mcm3m1f_cf_w_1_120_s_0_840=2.17e-11
.param mcm3m1f_ca_w_1_120_s_1_540=5.87e-05
.param mcm3m1f_cc_w_1_120_s_1_540=1.43e-11
.param mcm3m1f_cf_w_1_120_s_1_540=3.33e-11
.param mcm3m1f_ca_w_1_120_s_3_500=5.87e-05
.param mcm3m1f_cc_w_1_120_s_3_500=1.61e-12
.param mcm3m1f_cf_w_1_120_s_3_500=4.41e-11
.param mcm3m1d_ca_w_0_140_s_0_140=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_140=9.98e-11
.param mcm3m1d_cf_w_0_140_s_0_140=4.57e-12
.param mcm3m1d_ca_w_0_140_s_0_175=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_175=9.81e-11
.param mcm3m1d_cf_w_0_140_s_0_175=5.69e-12
.param mcm3m1d_ca_w_0_140_s_0_210=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_210=9.26e-11
.param mcm3m1d_cf_w_0_140_s_0_210=6.82e-12
.param mcm3m1d_ca_w_0_140_s_0_280=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_280=8.03e-11
.param mcm3m1d_cf_w_0_140_s_0_280=9.01e-12
.param mcm3m1d_ca_w_0_140_s_0_350=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_350=6.89e-11
.param mcm3m1d_cf_w_0_140_s_0_350=1.12e-11
.param mcm3m1d_ca_w_0_140_s_0_420=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_420=5.84e-11
.param mcm3m1d_cf_w_0_140_s_0_420=1.33e-11
.param mcm3m1d_ca_w_0_140_s_0_560=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_560=4.41e-11
.param mcm3m1d_cf_w_0_140_s_0_560=1.72e-11
.param mcm3m1d_ca_w_0_140_s_0_840=6.65e-05
.param mcm3m1d_cc_w_0_140_s_0_840=2.81e-11
.param mcm3m1d_cf_w_0_140_s_0_840=2.40e-11
.param mcm3m1d_ca_w_0_140_s_1_540=6.65e-05
.param mcm3m1d_cc_w_0_140_s_1_540=1.07e-11
.param mcm3m1d_cf_w_0_140_s_1_540=3.53e-11
.param mcm3m1d_ca_w_0_140_s_3_500=6.65e-05
.param mcm3m1d_cc_w_0_140_s_3_500=9.30e-13
.param mcm3m1d_cf_w_0_140_s_3_500=4.43e-11
.param mcm3m1d_ca_w_1_120_s_0_140=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_140=1.15e-10
.param mcm3m1d_cf_w_1_120_s_0_140=4.62e-12
.param mcm3m1d_ca_w_1_120_s_0_175=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_175=1.11e-10
.param mcm3m1d_cf_w_1_120_s_0_175=5.75e-12
.param mcm3m1d_ca_w_1_120_s_0_210=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_210=1.03e-10
.param mcm3m1d_cf_w_1_120_s_0_210=6.88e-12
.param mcm3m1d_ca_w_1_120_s_0_280=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_280=8.87e-11
.param mcm3m1d_cf_w_1_120_s_0_280=9.07e-12
.param mcm3m1d_ca_w_1_120_s_0_350=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_350=7.63e-11
.param mcm3m1d_cf_w_1_120_s_0_350=1.13e-11
.param mcm3m1d_ca_w_1_120_s_0_420=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_420=6.51e-11
.param mcm3m1d_cf_w_1_120_s_0_420=1.33e-11
.param mcm3m1d_ca_w_1_120_s_0_560=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_560=4.92e-11
.param mcm3m1d_cf_w_1_120_s_0_560=1.73e-11
.param mcm3m1d_ca_w_1_120_s_0_840=6.65e-05
.param mcm3m1d_cc_w_1_120_s_0_840=3.11e-11
.param mcm3m1d_cf_w_1_120_s_0_840=2.43e-11
.param mcm3m1d_ca_w_1_120_s_1_540=6.65e-05
.param mcm3m1d_cc_w_1_120_s_1_540=1.20e-11
.param mcm3m1d_cf_w_1_120_s_1_540=3.64e-11
.param mcm3m1d_ca_w_1_120_s_3_500=6.65e-05
.param mcm3m1d_cc_w_1_120_s_3_500=1.08e-12
.param mcm3m1d_cf_w_1_120_s_3_500=4.62e-11
.param mcm3m1p1_ca_w_0_140_s_0_140=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_140=9.86e-11
.param mcm3m1p1_cf_w_0_140_s_0_140=5.34e-12
.param mcm3m1p1_ca_w_0_140_s_0_175=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_175=9.67e-11
.param mcm3m1p1_cf_w_0_140_s_0_175=6.66e-12
.param mcm3m1p1_ca_w_0_140_s_0_210=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_210=9.06e-11
.param mcm3m1p1_cf_w_0_140_s_0_210=7.99e-12
.param mcm3m1p1_ca_w_0_140_s_0_280=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_280=7.85e-11
.param mcm3m1p1_cf_w_0_140_s_0_280=1.05e-11
.param mcm3m1p1_ca_w_0_140_s_0_350=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_350=6.65e-11
.param mcm3m1p1_cf_w_0_140_s_0_350=1.30e-11
.param mcm3m1p1_ca_w_0_140_s_0_420=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_420=5.61e-11
.param mcm3m1p1_cf_w_0_140_s_0_420=1.54e-11
.param mcm3m1p1_ca_w_0_140_s_0_560=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_560=4.20e-11
.param mcm3m1p1_cf_w_0_140_s_0_560=1.99e-11
.param mcm3m1p1_ca_w_0_140_s_0_840=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_0_840=2.56e-11
.param mcm3m1p1_cf_w_0_140_s_0_840=2.75e-11
.param mcm3m1p1_ca_w_0_140_s_1_540=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_1_540=8.79e-12
.param mcm3m1p1_cf_w_0_140_s_1_540=3.93e-11
.param mcm3m1p1_ca_w_0_140_s_3_500=7.78e-05
.param mcm3m1p1_cc_w_0_140_s_3_500=5.90e-13
.param mcm3m1p1_cf_w_0_140_s_3_500=4.72e-11
.param mcm3m1p1_ca_w_1_120_s_0_140=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_140=1.10e-10
.param mcm3m1p1_cf_w_1_120_s_0_140=5.45e-12
.param mcm3m1p1_ca_w_1_120_s_0_175=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_175=1.07e-10
.param mcm3m1p1_cf_w_1_120_s_0_175=6.77e-12
.param mcm3m1p1_ca_w_1_120_s_0_210=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_210=9.98e-11
.param mcm3m1p1_cf_w_1_120_s_0_210=8.09e-12
.param mcm3m1p1_ca_w_1_120_s_0_280=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_280=8.54e-11
.param mcm3m1p1_cf_w_1_120_s_0_280=1.06e-11
.param mcm3m1p1_ca_w_1_120_s_0_350=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_350=7.26e-11
.param mcm3m1p1_cf_w_1_120_s_0_350=1.32e-11
.param mcm3m1p1_ca_w_1_120_s_0_420=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_420=6.14e-11
.param mcm3m1p1_cf_w_1_120_s_0_420=1.56e-11
.param mcm3m1p1_ca_w_1_120_s_0_560=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_560=4.58e-11
.param mcm3m1p1_cf_w_1_120_s_0_560=2.01e-11
.param mcm3m1p1_ca_w_1_120_s_0_840=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_0_840=2.81e-11
.param mcm3m1p1_cf_w_1_120_s_0_840=2.79e-11
.param mcm3m1p1_ca_w_1_120_s_1_540=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_1_540=9.77e-12
.param mcm3m1p1_cf_w_1_120_s_1_540=4.05e-11
.param mcm3m1p1_ca_w_1_120_s_3_500=7.78e-05
.param mcm3m1p1_cc_w_1_120_s_3_500=6.25e-13
.param mcm3m1p1_cf_w_1_120_s_3_500=4.89e-11
.param mcm3m1l1_ca_w_0_140_s_0_140=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_140=9.23e-11
.param mcm3m1l1_cf_w_0_140_s_0_140=9.69e-12
.param mcm3m1l1_ca_w_0_140_s_0_175=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_175=8.99e-11
.param mcm3m1l1_cf_w_0_140_s_0_175=1.22e-11
.param mcm3m1l1_ca_w_0_140_s_0_210=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_210=8.35e-11
.param mcm3m1l1_cf_w_0_140_s_0_210=1.46e-11
.param mcm3m1l1_ca_w_0_140_s_0_280=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_280=7.03e-11
.param mcm3m1l1_cf_w_0_140_s_0_280=1.92e-11
.param mcm3m1l1_ca_w_0_140_s_0_350=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_350=5.81e-11
.param mcm3m1l1_cf_w_0_140_s_0_350=2.36e-11
.param mcm3m1l1_ca_w_0_140_s_0_420=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_420=4.76e-11
.param mcm3m1l1_cf_w_0_140_s_0_420=2.76e-11
.param mcm3m1l1_ca_w_0_140_s_0_560=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_560=3.32e-11
.param mcm3m1l1_cf_w_0_140_s_0_560=3.45e-11
.param mcm3m1l1_ca_w_0_140_s_0_840=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_0_840=1.76e-11
.param mcm3m1l1_cf_w_0_140_s_0_840=4.47e-11
.param mcm3m1l1_ca_w_0_140_s_1_540=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_1_540=4.42e-12
.param mcm3m1l1_cf_w_0_140_s_1_540=5.63e-11
.param mcm3m1l1_ca_w_0_140_s_3_500=1.47e-04
.param mcm3m1l1_cc_w_0_140_s_3_500=2.10e-13
.param mcm3m1l1_cf_w_0_140_s_3_500=6.09e-11
.param mcm3m1l1_ca_w_1_120_s_0_140=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_140=9.93e-11
.param mcm3m1l1_cf_w_1_120_s_0_140=9.78e-12
.param mcm3m1l1_ca_w_1_120_s_0_175=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_175=9.67e-11
.param mcm3m1l1_cf_w_1_120_s_0_175=1.23e-11
.param mcm3m1l1_ca_w_1_120_s_0_210=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_210=8.96e-11
.param mcm3m1l1_cf_w_1_120_s_0_210=1.47e-11
.param mcm3m1l1_ca_w_1_120_s_0_280=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_280=7.50e-11
.param mcm3m1l1_cf_w_1_120_s_0_280=1.93e-11
.param mcm3m1l1_ca_w_1_120_s_0_350=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_350=6.21e-11
.param mcm3m1l1_cf_w_1_120_s_0_350=2.36e-11
.param mcm3m1l1_ca_w_1_120_s_0_420=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_420=5.11e-11
.param mcm3m1l1_cf_w_1_120_s_0_420=2.76e-11
.param mcm3m1l1_ca_w_1_120_s_0_560=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_560=3.58e-11
.param mcm3m1l1_cf_w_1_120_s_0_560=3.47e-11
.param mcm3m1l1_ca_w_1_120_s_0_840=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_0_840=1.93e-11
.param mcm3m1l1_cf_w_1_120_s_0_840=4.52e-11
.param mcm3m1l1_ca_w_1_120_s_1_540=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_1_540=4.97e-12
.param mcm3m1l1_cf_w_1_120_s_1_540=5.75e-11
.param mcm3m1l1_ca_w_1_120_s_3_500=1.47e-04
.param mcm3m1l1_cc_w_1_120_s_3_500=2.35e-13
.param mcm3m1l1_cf_w_1_120_s_3_500=6.25e-11
.param mcm4m1f_ca_w_0_140_s_0_140=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_140=1.04e-10
.param mcm4m1f_cf_w_0_140_s_0_140=2.84e-12
.param mcm4m1f_ca_w_0_140_s_0_175=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_175=1.02e-10
.param mcm4m1f_cf_w_0_140_s_0_175=3.54e-12
.param mcm4m1f_ca_w_0_140_s_0_210=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_210=9.63e-11
.param mcm4m1f_cf_w_0_140_s_0_210=4.25e-12
.param mcm4m1f_ca_w_0_140_s_0_280=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_280=8.48e-11
.param mcm4m1f_cf_w_0_140_s_0_280=5.64e-12
.param mcm4m1f_ca_w_0_140_s_0_350=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_350=7.33e-11
.param mcm4m1f_cf_w_0_140_s_0_350=7.00e-12
.param mcm4m1f_ca_w_0_140_s_0_420=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_420=6.36e-11
.param mcm4m1f_cf_w_0_140_s_0_420=8.39e-12
.param mcm4m1f_ca_w_0_140_s_0_560=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_560=5.03e-11
.param mcm4m1f_cf_w_0_140_s_0_560=1.10e-11
.param mcm4m1f_ca_w_0_140_s_0_840=4.09e-05
.param mcm4m1f_cc_w_0_140_s_0_840=3.51e-11
.param mcm4m1f_cf_w_0_140_s_0_840=1.57e-11
.param mcm4m1f_ca_w_0_140_s_1_540=4.09e-05
.param mcm4m1f_cc_w_0_140_s_1_540=1.74e-11
.param mcm4m1f_cf_w_0_140_s_1_540=2.48e-11
.param mcm4m1f_ca_w_0_140_s_3_500=4.09e-05
.param mcm4m1f_cc_w_0_140_s_3_500=3.40e-12
.param mcm4m1f_cf_w_0_140_s_3_500=3.59e-11
.param mcm4m1f_ca_w_1_120_s_0_140=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_140=1.23e-10
.param mcm4m1f_cf_w_1_120_s_0_140=2.88e-12
.param mcm4m1f_ca_w_1_120_s_0_175=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_175=1.20e-10
.param mcm4m1f_cf_w_1_120_s_0_175=3.58e-12
.param mcm4m1f_ca_w_1_120_s_0_210=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_210=1.13e-10
.param mcm4m1f_cf_w_1_120_s_0_210=4.29e-12
.param mcm4m1f_ca_w_1_120_s_0_280=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_280=9.88e-11
.param mcm4m1f_cf_w_1_120_s_0_280=5.68e-12
.param mcm4m1f_ca_w_1_120_s_0_350=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_350=8.60e-11
.param mcm4m1f_cf_w_1_120_s_0_350=7.06e-12
.param mcm4m1f_ca_w_1_120_s_0_420=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_420=7.51e-11
.param mcm4m1f_cf_w_1_120_s_0_420=8.40e-12
.param mcm4m1f_ca_w_1_120_s_0_560=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_560=5.93e-11
.param mcm4m1f_cf_w_1_120_s_0_560=1.10e-11
.param mcm4m1f_ca_w_1_120_s_0_840=4.09e-05
.param mcm4m1f_cc_w_1_120_s_0_840=4.12e-11
.param mcm4m1f_cf_w_1_120_s_0_840=1.59e-11
.param mcm4m1f_ca_w_1_120_s_1_540=4.09e-05
.param mcm4m1f_cc_w_1_120_s_1_540=2.07e-11
.param mcm4m1f_cf_w_1_120_s_1_540=2.56e-11
.param mcm4m1f_ca_w_1_120_s_3_500=4.09e-05
.param mcm4m1f_cc_w_1_120_s_3_500=4.21e-12
.param mcm4m1f_cf_w_1_120_s_3_500=3.82e-11
.param mcm4m1d_ca_w_0_140_s_0_140=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_140=1.03e-10
.param mcm4m1d_cf_w_0_140_s_0_140=3.37e-12
.param mcm4m1d_ca_w_0_140_s_0_175=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_175=1.00e-10
.param mcm4m1d_cf_w_0_140_s_0_175=4.21e-12
.param mcm4m1d_ca_w_0_140_s_0_210=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_210=9.52e-11
.param mcm4m1d_cf_w_0_140_s_0_210=5.06e-12
.param mcm4m1d_ca_w_0_140_s_0_280=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_280=8.35e-11
.param mcm4m1d_cf_w_0_140_s_0_280=6.70e-12
.param mcm4m1d_ca_w_0_140_s_0_350=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_350=7.19e-11
.param mcm4m1d_cf_w_0_140_s_0_350=8.31e-12
.param mcm4m1d_ca_w_0_140_s_0_420=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_420=6.21e-11
.param mcm4m1d_cf_w_0_140_s_0_420=9.94e-12
.param mcm4m1d_ca_w_0_140_s_0_560=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_560=4.83e-11
.param mcm4m1d_cf_w_0_140_s_0_560=1.29e-11
.param mcm4m1d_ca_w_0_140_s_0_840=4.87e-05
.param mcm4m1d_cc_w_0_140_s_0_840=3.29e-11
.param mcm4m1d_cf_w_0_140_s_0_840=1.83e-11
.param mcm4m1d_ca_w_0_140_s_1_540=4.87e-05
.param mcm4m1d_cc_w_0_140_s_1_540=1.53e-11
.param mcm4m1d_cf_w_0_140_s_1_540=2.83e-11
.param mcm4m1d_ca_w_0_140_s_3_500=4.87e-05
.param mcm4m1d_cc_w_0_140_s_3_500=2.56e-12
.param mcm4m1d_cf_w_0_140_s_3_500=3.90e-11
.param mcm4m1d_ca_w_1_120_s_0_140=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_140=1.20e-10
.param mcm4m1d_cf_w_1_120_s_0_140=3.44e-12
.param mcm4m1d_ca_w_1_120_s_0_175=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_175=1.17e-10
.param mcm4m1d_cf_w_1_120_s_0_175=4.28e-12
.param mcm4m1d_ca_w_1_120_s_0_210=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_210=1.10e-10
.param mcm4m1d_cf_w_1_120_s_0_210=5.12e-12
.param mcm4m1d_ca_w_1_120_s_0_280=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_280=9.59e-11
.param mcm4m1d_cf_w_1_120_s_0_280=6.77e-12
.param mcm4m1d_ca_w_1_120_s_0_350=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_350=8.32e-11
.param mcm4m1d_cf_w_1_120_s_0_350=8.39e-12
.param mcm4m1d_ca_w_1_120_s_0_420=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_420=7.20e-11
.param mcm4m1d_cf_w_1_120_s_0_420=9.98e-12
.param mcm4m1d_ca_w_1_120_s_0_560=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_560=5.66e-11
.param mcm4m1d_cf_w_1_120_s_0_560=1.30e-11
.param mcm4m1d_ca_w_1_120_s_0_840=4.87e-05
.param mcm4m1d_cc_w_1_120_s_0_840=3.84e-11
.param mcm4m1d_cf_w_1_120_s_0_840=1.86e-11
.param mcm4m1d_ca_w_1_120_s_1_540=4.87e-05
.param mcm4m1d_cc_w_1_120_s_1_540=1.83e-11
.param mcm4m1d_cf_w_1_120_s_1_540=2.92e-11
.param mcm4m1d_ca_w_1_120_s_3_500=4.87e-05
.param mcm4m1d_cc_w_1_120_s_3_500=3.17e-12
.param mcm4m1d_cf_w_1_120_s_3_500=4.14e-11
.param mcm4m1p1_ca_w_0_140_s_0_140=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_140=1.02e-10
.param mcm4m1p1_cf_w_0_140_s_0_140=4.15e-12
.param mcm4m1p1_ca_w_0_140_s_0_175=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_175=9.91e-11
.param mcm4m1p1_cf_w_0_140_s_0_175=5.18e-12
.param mcm4m1p1_ca_w_0_140_s_0_210=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_210=9.32e-11
.param mcm4m1p1_cf_w_0_140_s_0_210=6.23e-12
.param mcm4m1p1_ca_w_0_140_s_0_280=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_280=8.17e-11
.param mcm4m1p1_cf_w_0_140_s_0_280=8.23e-12
.param mcm4m1p1_ca_w_0_140_s_0_350=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_350=6.97e-11
.param mcm4m1p1_cf_w_0_140_s_0_350=1.02e-11
.param mcm4m1p1_ca_w_0_140_s_0_420=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_420=6.00e-11
.param mcm4m1p1_cf_w_0_140_s_0_420=1.21e-11
.param mcm4m1p1_ca_w_0_140_s_0_560=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_560=4.62e-11
.param mcm4m1p1_cf_w_0_140_s_0_560=1.57e-11
.param mcm4m1p1_ca_w_0_140_s_0_840=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_0_840=3.03e-11
.param mcm4m1p1_cf_w_0_140_s_0_840=2.20e-11
.param mcm4m1p1_ca_w_0_140_s_1_540=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_1_540=1.31e-11
.param mcm4m1p1_cf_w_0_140_s_1_540=3.28e-11
.param mcm4m1p1_ca_w_0_140_s_3_500=6.00e-05
.param mcm4m1p1_cc_w_0_140_s_3_500=1.84e-12
.param mcm4m1p1_cf_w_0_140_s_3_500=4.27e-11
.param mcm4m1p1_ca_w_1_120_s_0_140=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_140=1.17e-10
.param mcm4m1p1_cf_w_1_120_s_0_140=4.31e-12
.param mcm4m1p1_ca_w_1_120_s_0_175=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_175=1.13e-10
.param mcm4m1p1_cf_w_1_120_s_0_175=5.32e-12
.param mcm4m1p1_ca_w_1_120_s_0_210=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_210=1.07e-10
.param mcm4m1p1_cf_w_1_120_s_0_210=6.34e-12
.param mcm4m1p1_ca_w_1_120_s_0_280=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_280=9.24e-11
.param mcm4m1p1_cf_w_1_120_s_0_280=8.35e-12
.param mcm4m1p1_ca_w_1_120_s_0_350=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_350=7.96e-11
.param mcm4m1p1_cf_w_1_120_s_0_350=1.03e-11
.param mcm4m1p1_ca_w_1_120_s_0_420=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_420=6.88e-11
.param mcm4m1p1_cf_w_1_120_s_0_420=1.22e-11
.param mcm4m1p1_ca_w_1_120_s_0_560=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_560=5.30e-11
.param mcm4m1p1_cf_w_1_120_s_0_560=1.59e-11
.param mcm4m1p1_ca_w_1_120_s_0_840=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_0_840=3.52e-11
.param mcm4m1p1_cf_w_1_120_s_0_840=2.23e-11
.param mcm4m1p1_ca_w_1_120_s_1_540=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_1_540=1.57e-11
.param mcm4m1p1_cf_w_1_120_s_1_540=3.38e-11
.param mcm4m1p1_ca_w_1_120_s_3_500=6.00e-05
.param mcm4m1p1_cc_w_1_120_s_3_500=2.33e-12
.param mcm4m1p1_cf_w_1_120_s_3_500=4.52e-11
.param mcm4m1l1_ca_w_0_140_s_0_140=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_140=9.48e-11
.param mcm4m1l1_cf_w_0_140_s_0_140=8.49e-12
.param mcm4m1l1_ca_w_0_140_s_0_175=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_175=9.24e-11
.param mcm4m1l1_cf_w_0_140_s_0_175=1.07e-11
.param mcm4m1l1_ca_w_0_140_s_0_210=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_210=8.59e-11
.param mcm4m1l1_cf_w_0_140_s_0_210=1.29e-11
.param mcm4m1l1_ca_w_0_140_s_0_280=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_280=7.35e-11
.param mcm4m1l1_cf_w_0_140_s_0_280=1.69e-11
.param mcm4m1l1_ca_w_0_140_s_0_350=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_350=6.15e-11
.param mcm4m1l1_cf_w_0_140_s_0_350=2.07e-11
.param mcm4m1l1_ca_w_0_140_s_0_420=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_420=5.10e-11
.param mcm4m1l1_cf_w_0_140_s_0_420=2.42e-11
.param mcm4m1l1_ca_w_0_140_s_0_560=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_560=3.72e-11
.param mcm4m1l1_cf_w_0_140_s_0_560=3.04e-11
.param mcm4m1l1_ca_w_0_140_s_0_840=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_0_840=2.20e-11
.param mcm4m1l1_cf_w_0_140_s_0_840=3.97e-11
.param mcm4m1l1_ca_w_0_140_s_1_540=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_1_540=7.54e-12
.param mcm4m1l1_cf_w_0_140_s_1_540=5.16e-11
.param mcm4m1l1_ca_w_0_140_s_3_500=1.29e-04
.param mcm4m1l1_cc_w_0_140_s_3_500=7.50e-13
.param mcm4m1l1_cf_w_0_140_s_3_500=5.84e-11
.param mcm4m1l1_ca_w_1_120_s_0_140=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_140=1.06e-10
.param mcm4m1l1_cf_w_1_120_s_0_140=8.63e-12
.param mcm4m1l1_ca_w_1_120_s_0_175=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_175=1.03e-10
.param mcm4m1l1_cf_w_1_120_s_0_175=1.08e-11
.param mcm4m1l1_ca_w_1_120_s_0_210=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_210=9.61e-11
.param mcm4m1l1_cf_w_1_120_s_0_210=1.30e-11
.param mcm4m1l1_ca_w_1_120_s_0_280=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_280=8.18e-11
.param mcm4m1l1_cf_w_1_120_s_0_280=1.70e-11
.param mcm4m1l1_ca_w_1_120_s_0_350=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_350=6.92e-11
.param mcm4m1l1_cf_w_1_120_s_0_350=2.08e-11
.param mcm4m1l1_ca_w_1_120_s_0_420=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_420=5.81e-11
.param mcm4m1l1_cf_w_1_120_s_0_420=2.43e-11
.param mcm4m1l1_ca_w_1_120_s_0_560=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_560=4.30e-11
.param mcm4m1l1_cf_w_1_120_s_0_560=3.05e-11
.param mcm4m1l1_ca_w_1_120_s_0_840=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_0_840=2.62e-11
.param mcm4m1l1_cf_w_1_120_s_0_840=4.01e-11
.param mcm4m1l1_ca_w_1_120_s_1_540=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_1_540=9.81e-12
.param mcm4m1l1_cf_w_1_120_s_1_540=5.30e-11
.param mcm4m1l1_ca_w_1_120_s_3_500=1.29e-04
.param mcm4m1l1_cc_w_1_120_s_3_500=1.05e-12
.param mcm4m1l1_cf_w_1_120_s_3_500=6.13e-11
.param mcm5m1f_ca_w_0_140_s_0_140=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_140=1.04e-10
.param mcm5m1f_cf_w_0_140_s_0_140=2.45e-12
.param mcm5m1f_ca_w_0_140_s_0_175=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_175=1.02e-10
.param mcm5m1f_cf_w_0_140_s_0_175=3.06e-12
.param mcm5m1f_ca_w_0_140_s_0_210=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_210=9.71e-11
.param mcm5m1f_cf_w_0_140_s_0_210=3.68e-12
.param mcm5m1f_ca_w_0_140_s_0_280=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_280=8.58e-11
.param mcm5m1f_cf_w_0_140_s_0_280=4.88e-12
.param mcm5m1f_ca_w_0_140_s_0_350=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_350=7.46e-11
.param mcm5m1f_cf_w_0_140_s_0_350=6.06e-12
.param mcm5m1f_ca_w_0_140_s_0_420=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_420=6.50e-11
.param mcm5m1f_cf_w_0_140_s_0_420=7.28e-12
.param mcm5m1f_ca_w_0_140_s_0_560=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_560=5.17e-11
.param mcm5m1f_cf_w_0_140_s_0_560=9.53e-12
.param mcm5m1f_ca_w_0_140_s_0_840=3.53e-05
.param mcm5m1f_cc_w_0_140_s_0_840=3.70e-11
.param mcm5m1f_cf_w_0_140_s_0_840=1.37e-11
.param mcm5m1f_ca_w_0_140_s_1_540=3.53e-05
.param mcm5m1f_cc_w_0_140_s_1_540=1.97e-11
.param mcm5m1f_cf_w_0_140_s_1_540=2.20e-11
.param mcm5m1f_ca_w_0_140_s_3_500=3.53e-05
.param mcm5m1f_cc_w_0_140_s_3_500=4.95e-12
.param mcm5m1f_cf_w_0_140_s_3_500=3.32e-11
.param mcm5m1f_ca_w_1_120_s_0_140=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_140=1.25e-10
.param mcm5m1f_cf_w_1_120_s_0_140=2.49e-12
.param mcm5m1f_ca_w_1_120_s_0_175=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_175=1.23e-10
.param mcm5m1f_cf_w_1_120_s_0_175=3.10e-12
.param mcm5m1f_ca_w_1_120_s_0_210=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_210=1.16e-10
.param mcm5m1f_cf_w_1_120_s_0_210=3.72e-12
.param mcm5m1f_ca_w_1_120_s_0_280=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_280=1.02e-10
.param mcm5m1f_cf_w_1_120_s_0_280=4.92e-12
.param mcm5m1f_ca_w_1_120_s_0_350=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_350=8.91e-11
.param mcm5m1f_cf_w_1_120_s_0_350=6.11e-12
.param mcm5m1f_ca_w_1_120_s_0_420=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_420=7.82e-11
.param mcm5m1f_cf_w_1_120_s_0_420=7.29e-12
.param mcm5m1f_ca_w_1_120_s_0_560=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_560=6.26e-11
.param mcm5m1f_cf_w_1_120_s_0_560=9.56e-12
.param mcm5m1f_ca_w_1_120_s_0_840=3.53e-05
.param mcm5m1f_cc_w_1_120_s_0_840=4.47e-11
.param mcm5m1f_cf_w_1_120_s_0_840=1.38e-11
.param mcm5m1f_ca_w_1_120_s_1_540=3.53e-05
.param mcm5m1f_cc_w_1_120_s_1_540=2.43e-11
.param mcm5m1f_cf_w_1_120_s_1_540=2.26e-11
.param mcm5m1f_ca_w_1_120_s_3_500=3.53e-05
.param mcm5m1f_cc_w_1_120_s_3_500=6.46e-12
.param mcm5m1f_cf_w_1_120_s_3_500=3.55e-11
.param mcm5m1d_ca_w_0_140_s_0_140=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_140=1.03e-10
.param mcm5m1d_cf_w_0_140_s_0_140=2.99e-12
.param mcm5m1d_ca_w_0_140_s_0_175=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_175=1.01e-10
.param mcm5m1d_cf_w_0_140_s_0_175=3.73e-12
.param mcm5m1d_ca_w_0_140_s_0_210=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_210=9.56e-11
.param mcm5m1d_cf_w_0_140_s_0_210=4.49e-12
.param mcm5m1d_ca_w_0_140_s_0_280=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_280=8.45e-11
.param mcm5m1d_cf_w_0_140_s_0_280=5.95e-12
.param mcm5m1d_ca_w_0_140_s_0_350=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_350=7.26e-11
.param mcm5m1d_cf_w_0_140_s_0_350=7.38e-12
.param mcm5m1d_ca_w_0_140_s_0_420=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_420=6.30e-11
.param mcm5m1d_cf_w_0_140_s_0_420=8.82e-12
.param mcm5m1d_ca_w_0_140_s_0_560=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_560=5.00e-11
.param mcm5m1d_cf_w_0_140_s_0_560=1.15e-11
.param mcm5m1d_ca_w_0_140_s_0_840=4.31e-05
.param mcm5m1d_cc_w_0_140_s_0_840=3.48e-11
.param mcm5m1d_cf_w_0_140_s_0_840=1.64e-11
.param mcm5m1d_ca_w_0_140_s_1_540=4.31e-05
.param mcm5m1d_cc_w_0_140_s_1_540=1.75e-11
.param mcm5m1d_cf_w_0_140_s_1_540=2.56e-11
.param mcm5m1d_ca_w_0_140_s_3_500=4.31e-05
.param mcm5m1d_cc_w_0_140_s_3_500=3.87e-12
.param mcm5m1d_cf_w_0_140_s_3_500=3.66e-11
.param mcm5m1d_ca_w_1_120_s_0_140=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_140=1.23e-10
.param mcm5m1d_cf_w_1_120_s_0_140=3.06e-12
.param mcm5m1d_ca_w_1_120_s_0_175=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_175=1.20e-10
.param mcm5m1d_cf_w_1_120_s_0_175=3.80e-12
.param mcm5m1d_ca_w_1_120_s_0_210=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_210=1.13e-10
.param mcm5m1d_cf_w_1_120_s_0_210=4.55e-12
.param mcm5m1d_ca_w_1_120_s_0_280=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_280=9.88e-11
.param mcm5m1d_cf_w_1_120_s_0_280=6.01e-12
.param mcm5m1d_ca_w_1_120_s_0_350=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_350=8.63e-11
.param mcm5m1d_cf_w_1_120_s_0_350=7.45e-12
.param mcm5m1d_ca_w_1_120_s_0_420=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_420=7.51e-11
.param mcm5m1d_cf_w_1_120_s_0_420=8.86e-12
.param mcm5m1d_ca_w_1_120_s_0_560=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_560=5.97e-11
.param mcm5m1d_cf_w_1_120_s_0_560=1.16e-11
.param mcm5m1d_ca_w_1_120_s_0_840=4.31e-05
.param mcm5m1d_cc_w_1_120_s_0_840=4.17e-11
.param mcm5m1d_cf_w_1_120_s_0_840=1.66e-11
.param mcm5m1d_ca_w_1_120_s_1_540=4.31e-05
.param mcm5m1d_cc_w_1_120_s_1_540=2.17e-11
.param mcm5m1d_cf_w_1_120_s_1_540=2.63e-11
.param mcm5m1d_ca_w_1_120_s_3_500=4.31e-05
.param mcm5m1d_cc_w_1_120_s_3_500=5.18e-12
.param mcm5m1d_cf_w_1_120_s_3_500=3.92e-11
.param mcm5m1p1_ca_w_0_140_s_0_140=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_140=1.02e-10
.param mcm5m1p1_cf_w_0_140_s_0_140=3.77e-12
.param mcm5m1p1_ca_w_0_140_s_0_175=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_175=9.98e-11
.param mcm5m1p1_cf_w_0_140_s_0_175=4.71e-12
.param mcm5m1p1_ca_w_0_140_s_0_210=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_210=9.41e-11
.param mcm5m1p1_cf_w_0_140_s_0_210=5.65e-12
.param mcm5m1p1_ca_w_0_140_s_0_280=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_280=8.27e-11
.param mcm5m1p1_cf_w_0_140_s_0_280=7.48e-12
.param mcm5m1p1_ca_w_0_140_s_0_350=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_350=7.09e-11
.param mcm5m1p1_cf_w_0_140_s_0_350=9.24e-12
.param mcm5m1p1_ca_w_0_140_s_0_420=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_420=6.10e-11
.param mcm5m1p1_cf_w_0_140_s_0_420=1.10e-11
.param mcm5m1p1_ca_w_0_140_s_0_560=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_560=4.76e-11
.param mcm5m1p1_cf_w_0_140_s_0_560=1.43e-11
.param mcm5m1p1_ca_w_0_140_s_0_840=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_0_840=3.22e-11
.param mcm5m1p1_cf_w_0_140_s_0_840=2.01e-11
.param mcm5m1p1_ca_w_0_140_s_1_540=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_1_540=1.52e-11
.param mcm5m1p1_cf_w_0_140_s_1_540=3.03e-11
.param mcm5m1p1_ca_w_0_140_s_3_500=5.44e-05
.param mcm5m1p1_cc_w_0_140_s_3_500=2.95e-12
.param mcm5m1p1_cf_w_0_140_s_3_500=4.08e-11
.param mcm5m1p1_ca_w_1_120_s_0_140=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_140=1.20e-10
.param mcm5m1p1_cf_w_1_120_s_0_140=3.92e-12
.param mcm5m1p1_ca_w_1_120_s_0_175=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_175=1.16e-10
.param mcm5m1p1_cf_w_1_120_s_0_175=4.86e-12
.param mcm5m1p1_ca_w_1_120_s_0_210=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_210=1.10e-10
.param mcm5m1p1_cf_w_1_120_s_0_210=5.78e-12
.param mcm5m1p1_ca_w_1_120_s_0_280=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_280=9.54e-11
.param mcm5m1p1_cf_w_1_120_s_0_280=7.61e-12
.param mcm5m1p1_ca_w_1_120_s_0_350=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_350=8.27e-11
.param mcm5m1p1_cf_w_1_120_s_0_350=9.40e-12
.param mcm5m1p1_ca_w_1_120_s_0_420=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_420=7.19e-11
.param mcm5m1p1_cf_w_1_120_s_0_420=1.12e-11
.param mcm5m1p1_ca_w_1_120_s_0_560=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_560=5.62e-11
.param mcm5m1p1_cf_w_1_120_s_0_560=1.44e-11
.param mcm5m1p1_ca_w_1_120_s_0_840=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_0_840=3.86e-11
.param mcm5m1p1_cf_w_1_120_s_0_840=2.04e-11
.param mcm5m1p1_ca_w_1_120_s_1_540=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_1_540=1.91e-11
.param mcm5m1p1_cf_w_1_120_s_1_540=3.13e-11
.param mcm5m1p1_ca_w_1_120_s_3_500=5.44e-05
.param mcm5m1p1_cc_w_1_120_s_3_500=4.05e-12
.param mcm5m1p1_cf_w_1_120_s_3_500=4.36e-11
.param mcm5m1l1_ca_w_0_140_s_0_140=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_140=9.56e-11
.param mcm5m1l1_cf_w_0_140_s_0_140=8.10e-12
.param mcm5m1l1_ca_w_0_140_s_0_175=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_175=9.31e-11
.param mcm5m1l1_cf_w_0_140_s_0_175=1.02e-11
.param mcm5m1l1_ca_w_0_140_s_0_210=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_210=8.67e-11
.param mcm5m1l1_cf_w_0_140_s_0_210=1.23e-11
.param mcm5m1l1_ca_w_0_140_s_0_280=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_280=7.45e-11
.param mcm5m1l1_cf_w_0_140_s_0_280=1.62e-11
.param mcm5m1l1_ca_w_0_140_s_0_350=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_350=6.24e-11
.param mcm5m1l1_cf_w_0_140_s_0_350=1.97e-11
.param mcm5m1l1_ca_w_0_140_s_0_420=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_420=5.25e-11
.param mcm5m1l1_cf_w_0_140_s_0_420=2.31e-11
.param mcm5m1l1_ca_w_0_140_s_0_560=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_560=3.86e-11
.param mcm5m1l1_cf_w_0_140_s_0_560=2.90e-11
.param mcm5m1l1_ca_w_0_140_s_0_840=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_0_840=2.38e-11
.param mcm5m1l1_cf_w_0_140_s_0_840=3.80e-11
.param mcm5m1l1_ca_w_0_140_s_1_540=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_1_540=9.09e-12
.param mcm5m1l1_cf_w_0_140_s_1_540=4.98e-11
.param mcm5m1l1_ca_w_0_140_s_3_500=1.23e-04
.param mcm5m1l1_cc_w_0_140_s_3_500=1.36e-12
.param mcm5m1l1_cf_w_0_140_s_3_500=5.74e-11
.param mcm5m1l1_ca_w_1_120_s_0_140=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_140=1.09e-10
.param mcm5m1l1_cf_w_1_120_s_0_140=8.26e-12
.param mcm5m1l1_ca_w_1_120_s_0_175=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_175=1.06e-10
.param mcm5m1l1_cf_w_1_120_s_0_175=1.04e-11
.param mcm5m1l1_ca_w_1_120_s_0_210=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_210=9.89e-11
.param mcm5m1l1_cf_w_1_120_s_0_210=1.24e-11
.param mcm5m1l1_ca_w_1_120_s_0_280=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_280=8.49e-11
.param mcm5m1l1_cf_w_1_120_s_0_280=1.63e-11
.param mcm5m1l1_ca_w_1_120_s_0_350=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_350=7.23e-11
.param mcm5m1l1_cf_w_1_120_s_0_350=1.99e-11
.param mcm5m1l1_ca_w_1_120_s_0_420=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_420=6.11e-11
.param mcm5m1l1_cf_w_1_120_s_0_420=2.33e-11
.param mcm5m1l1_ca_w_1_120_s_0_560=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_560=4.62e-11
.param mcm5m1l1_cf_w_1_120_s_0_560=2.91e-11
.param mcm5m1l1_ca_w_1_120_s_0_840=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_0_840=2.95e-11
.param mcm5m1l1_cf_w_1_120_s_0_840=3.83e-11
.param mcm5m1l1_ca_w_1_120_s_1_540=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_1_540=1.26e-11
.param mcm5m1l1_cf_w_1_120_s_1_540=5.10e-11
.param mcm5m1l1_ca_w_1_120_s_3_500=1.23e-04
.param mcm5m1l1_cc_w_1_120_s_3_500=2.20e-12
.param mcm5m1l1_cf_w_1_120_s_3_500=6.09e-11
.param mcrdlm1f_ca_w_0_140_s_0_140=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_140=1.05e-10
.param mcrdlm1f_cf_w_0_140_s_0_140=2.00e-12
.param mcrdlm1f_ca_w_0_140_s_0_175=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_175=1.03e-10
.param mcrdlm1f_cf_w_0_140_s_0_175=2.49e-12
.param mcrdlm1f_ca_w_0_140_s_0_210=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_210=9.77e-11
.param mcrdlm1f_cf_w_0_140_s_0_210=3.00e-12
.param mcrdlm1f_ca_w_0_140_s_0_280=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_280=8.68e-11
.param mcrdlm1f_cf_w_0_140_s_0_280=3.98e-12
.param mcrdlm1f_ca_w_0_140_s_0_350=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_350=7.54e-11
.param mcrdlm1f_cf_w_0_140_s_0_350=4.94e-12
.param mcrdlm1f_ca_w_0_140_s_0_420=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_420=6.65e-11
.param mcrdlm1f_cf_w_0_140_s_0_420=5.94e-12
.param mcrdlm1f_ca_w_0_140_s_0_560=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_560=5.36e-11
.param mcrdlm1f_cf_w_0_140_s_0_560=7.76e-12
.param mcrdlm1f_ca_w_0_140_s_0_840=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_0_840=3.94e-11
.param mcrdlm1f_cf_w_0_140_s_0_840=1.12e-11
.param mcrdlm1f_ca_w_0_140_s_1_540=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_1_540=2.30e-11
.param mcrdlm1f_cf_w_0_140_s_1_540=1.83e-11
.param mcrdlm1f_ca_w_0_140_s_3_500=2.87e-05
.param mcrdlm1f_cc_w_0_140_s_3_500=8.05e-12
.param mcrdlm1f_cf_w_0_140_s_3_500=2.92e-11
.param mcrdlm1f_ca_w_1_120_s_0_140=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_140=1.29e-10
.param mcrdlm1f_cf_w_1_120_s_0_140=2.04e-12
.param mcrdlm1f_ca_w_1_120_s_0_175=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_175=1.25e-10
.param mcrdlm1f_cf_w_1_120_s_0_175=2.54e-12
.param mcrdlm1f_ca_w_1_120_s_0_210=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_210=1.19e-10
.param mcrdlm1f_cf_w_1_120_s_0_210=3.04e-12
.param mcrdlm1f_ca_w_1_120_s_0_280=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_280=1.05e-10
.param mcrdlm1f_cf_w_1_120_s_0_280=4.03e-12
.param mcrdlm1f_ca_w_1_120_s_0_350=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_350=9.30e-11
.param mcrdlm1f_cf_w_1_120_s_0_350=5.00e-12
.param mcrdlm1f_ca_w_1_120_s_0_420=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_420=8.20e-11
.param mcrdlm1f_cf_w_1_120_s_0_420=5.95e-12
.param mcrdlm1f_ca_w_1_120_s_0_560=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_560=6.69e-11
.param mcrdlm1f_cf_w_1_120_s_0_560=7.81e-12
.param mcrdlm1f_ca_w_1_120_s_0_840=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_0_840=4.96e-11
.param mcrdlm1f_cf_w_1_120_s_0_840=1.13e-11
.param mcrdlm1f_ca_w_1_120_s_1_540=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_1_540=2.99e-11
.param mcrdlm1f_cf_w_1_120_s_1_540=1.88e-11
.param mcrdlm1f_ca_w_1_120_s_3_500=2.87e-05
.param mcrdlm1f_cc_w_1_120_s_3_500=1.14e-11
.param mcrdlm1f_cf_w_1_120_s_3_500=3.12e-11
.param mcrdlm1d_ca_w_0_140_s_0_140=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_140=1.04e-10
.param mcrdlm1d_cf_w_0_140_s_0_140=2.53e-12
.param mcrdlm1d_ca_w_0_140_s_0_175=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_175=1.02e-10
.param mcrdlm1d_cf_w_0_140_s_0_175=3.16e-12
.param mcrdlm1d_ca_w_0_140_s_0_210=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_210=9.66e-11
.param mcrdlm1d_cf_w_0_140_s_0_210=3.80e-12
.param mcrdlm1d_ca_w_0_140_s_0_280=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_280=8.55e-11
.param mcrdlm1d_cf_w_0_140_s_0_280=5.04e-12
.param mcrdlm1d_ca_w_0_140_s_0_350=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_350=7.40e-11
.param mcrdlm1d_cf_w_0_140_s_0_350=6.25e-12
.param mcrdlm1d_ca_w_0_140_s_0_420=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_420=6.49e-11
.param mcrdlm1d_cf_w_0_140_s_0_420=7.49e-12
.param mcrdlm1d_ca_w_0_140_s_0_560=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_560=5.17e-11
.param mcrdlm1d_cf_w_0_140_s_0_560=9.74e-12
.param mcrdlm1d_ca_w_0_140_s_0_840=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_0_840=3.72e-11
.param mcrdlm1d_cf_w_0_140_s_0_840=1.39e-11
.param mcrdlm1d_ca_w_0_140_s_1_540=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_1_540=2.08e-11
.param mcrdlm1d_cf_w_0_140_s_1_540=2.22e-11
.param mcrdlm1d_ca_w_0_140_s_3_500=3.65e-05
.param mcrdlm1d_cc_w_0_140_s_3_500=6.54e-12
.param mcrdlm1d_cf_w_0_140_s_3_500=3.32e-11
.param mcrdlm1d_ca_w_1_120_s_0_140=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_140=1.26e-10
.param mcrdlm1d_cf_w_1_120_s_0_140=2.61e-12
.param mcrdlm1d_ca_w_1_120_s_0_175=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_175=1.23e-10
.param mcrdlm1d_cf_w_1_120_s_0_175=3.24e-12
.param mcrdlm1d_ca_w_1_120_s_0_210=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_210=1.16e-10
.param mcrdlm1d_cf_w_1_120_s_0_210=3.87e-12
.param mcrdlm1d_ca_w_1_120_s_0_280=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_280=1.03e-10
.param mcrdlm1d_cf_w_1_120_s_0_280=5.12e-12
.param mcrdlm1d_ca_w_1_120_s_0_350=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_350=9.03e-11
.param mcrdlm1d_cf_w_1_120_s_0_350=6.34e-12
.param mcrdlm1d_ca_w_1_120_s_0_420=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_420=7.95e-11
.param mcrdlm1d_cf_w_1_120_s_0_420=7.53e-12
.param mcrdlm1d_ca_w_1_120_s_0_560=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_560=6.41e-11
.param mcrdlm1d_cf_w_1_120_s_0_560=9.83e-12
.param mcrdlm1d_ca_w_1_120_s_0_840=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_0_840=4.68e-11
.param mcrdlm1d_cf_w_1_120_s_0_840=1.41e-11
.param mcrdlm1d_ca_w_1_120_s_1_540=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_1_540=2.72e-11
.param mcrdlm1d_cf_w_1_120_s_1_540=2.27e-11
.param mcrdlm1d_ca_w_1_120_s_3_500=3.65e-05
.param mcrdlm1d_cc_w_1_120_s_3_500=9.66e-12
.param mcrdlm1d_cf_w_1_120_s_3_500=3.56e-11
.param mcrdlm1p1_ca_w_0_140_s_0_140=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_140=1.03e-10
.param mcrdlm1p1_cf_w_0_140_s_0_140=3.31e-12
.param mcrdlm1p1_ca_w_0_140_s_0_175=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_175=1.01e-10
.param mcrdlm1p1_cf_w_0_140_s_0_175=4.13e-12
.param mcrdlm1p1_ca_w_0_140_s_0_210=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_210=9.50e-11
.param mcrdlm1p1_cf_w_0_140_s_0_210=4.96e-12
.param mcrdlm1p1_ca_w_0_140_s_0_280=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_280=8.37e-11
.param mcrdlm1p1_cf_w_0_140_s_0_280=6.57e-12
.param mcrdlm1p1_ca_w_0_140_s_0_350=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_350=7.21e-11
.param mcrdlm1p1_cf_w_0_140_s_0_350=8.13e-12
.param mcrdlm1p1_ca_w_0_140_s_0_420=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_420=6.25e-11
.param mcrdlm1p1_cf_w_0_140_s_0_420=9.69e-12
.param mcrdlm1p1_ca_w_0_140_s_0_560=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_560=4.94e-11
.param mcrdlm1p1_cf_w_0_140_s_0_560=1.25e-11
.param mcrdlm1p1_ca_w_0_140_s_0_840=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_0_840=3.47e-11
.param mcrdlm1p1_cf_w_0_140_s_0_840=1.77e-11
.param mcrdlm1p1_ca_w_0_140_s_1_540=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_1_540=1.81e-11
.param mcrdlm1p1_cf_w_0_140_s_1_540=2.71e-11
.param mcrdlm1p1_ca_w_0_140_s_3_500=4.78e-05
.param mcrdlm1p1_cc_w_0_140_s_3_500=5.22e-12
.param mcrdlm1p1_cf_w_0_140_s_3_500=3.80e-11
.param mcrdlm1p1_ca_w_1_120_s_0_140=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_140=1.23e-10
.param mcrdlm1p1_cf_w_1_120_s_0_140=3.46e-12
.param mcrdlm1p1_ca_w_1_120_s_0_175=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_175=1.20e-10
.param mcrdlm1p1_cf_w_1_120_s_0_175=4.29e-12
.param mcrdlm1p1_ca_w_1_120_s_0_210=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_210=1.13e-10
.param mcrdlm1p1_cf_w_1_120_s_0_210=5.11e-12
.param mcrdlm1p1_ca_w_1_120_s_0_280=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_280=9.92e-11
.param mcrdlm1p1_cf_w_1_120_s_0_280=6.72e-12
.param mcrdlm1p1_ca_w_1_120_s_0_350=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_350=8.63e-11
.param mcrdlm1p1_cf_w_1_120_s_0_350=8.28e-12
.param mcrdlm1p1_ca_w_1_120_s_0_420=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_420=7.59e-11
.param mcrdlm1p1_cf_w_1_120_s_0_420=9.81e-12
.param mcrdlm1p1_ca_w_1_120_s_0_560=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_560=6.08e-11
.param mcrdlm1p1_cf_w_1_120_s_0_560=1.27e-11
.param mcrdlm1p1_ca_w_1_120_s_0_840=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_0_840=4.35e-11
.param mcrdlm1p1_cf_w_1_120_s_0_840=1.79e-11
.param mcrdlm1p1_ca_w_1_120_s_1_540=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_1_540=2.44e-11
.param mcrdlm1p1_cf_w_1_120_s_1_540=2.79e-11
.param mcrdlm1p1_ca_w_1_120_s_3_500=4.78e-05
.param mcrdlm1p1_cc_w_1_120_s_3_500=8.04e-12
.param mcrdlm1p1_cf_w_1_120_s_3_500=4.07e-11
.param mcrdlm1l1_ca_w_0_140_s_0_140=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_140=9.58e-11
.param mcrdlm1l1_cf_w_0_140_s_0_140=7.64e-12
.param mcrdlm1l1_ca_w_0_140_s_0_175=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_175=9.30e-11
.param mcrdlm1l1_cf_w_0_140_s_0_175=9.66e-12
.param mcrdlm1l1_ca_w_0_140_s_0_210=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_210=8.74e-11
.param mcrdlm1l1_cf_w_0_140_s_0_210=1.16e-11
.param mcrdlm1l1_ca_w_0_140_s_0_280=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_280=7.52e-11
.param mcrdlm1l1_cf_w_0_140_s_0_280=1.53e-11
.param mcrdlm1l1_ca_w_0_140_s_0_350=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_350=6.40e-11
.param mcrdlm1l1_cf_w_0_140_s_0_350=1.86e-11
.param mcrdlm1l1_ca_w_0_140_s_0_420=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_420=5.38e-11
.param mcrdlm1l1_cf_w_0_140_s_0_420=2.18e-11
.param mcrdlm1l1_ca_w_0_140_s_0_560=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_560=4.04e-11
.param mcrdlm1l1_cf_w_0_140_s_0_560=2.73e-11
.param mcrdlm1l1_ca_w_0_140_s_0_840=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_0_840=2.60e-11
.param mcrdlm1l1_cf_w_0_140_s_0_840=3.58e-11
.param mcrdlm1l1_ca_w_0_140_s_1_540=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_1_540=1.14e-11
.param mcrdlm1l1_cf_w_0_140_s_1_540=4.74e-11
.param mcrdlm1l1_ca_w_0_140_s_3_500=1.17e-04
.param mcrdlm1l1_cc_w_0_140_s_3_500=2.65e-12
.param mcrdlm1l1_cf_w_0_140_s_3_500=5.60e-11
.param mcrdlm1l1_ca_w_1_120_s_0_140=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_140=1.12e-10
.param mcrdlm1l1_cf_w_1_120_s_0_140=7.79e-12
.param mcrdlm1l1_ca_w_1_120_s_0_175=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_175=1.09e-10
.param mcrdlm1l1_cf_w_1_120_s_0_175=9.81e-12
.param mcrdlm1l1_ca_w_1_120_s_0_210=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_210=1.03e-10
.param mcrdlm1l1_cf_w_1_120_s_0_210=1.17e-11
.param mcrdlm1l1_ca_w_1_120_s_0_280=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_280=8.88e-11
.param mcrdlm1l1_cf_w_1_120_s_0_280=1.54e-11
.param mcrdlm1l1_ca_w_1_120_s_0_350=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_350=7.58e-11
.param mcrdlm1l1_cf_w_1_120_s_0_350=1.88e-11
.param mcrdlm1l1_ca_w_1_120_s_0_420=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_420=6.55e-11
.param mcrdlm1l1_cf_w_1_120_s_0_420=2.19e-11
.param mcrdlm1l1_ca_w_1_120_s_0_560=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_560=5.06e-11
.param mcrdlm1l1_cf_w_1_120_s_0_560=2.74e-11
.param mcrdlm1l1_ca_w_1_120_s_0_840=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_0_840=3.41e-11
.param mcrdlm1l1_cf_w_1_120_s_0_840=3.61e-11
.param mcrdlm1l1_ca_w_1_120_s_1_540=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_1_540=1.72e-11
.param mcrdlm1l1_cf_w_1_120_s_1_540=4.86e-11
.param mcrdlm1l1_ca_w_1_120_s_3_500=1.17e-04
.param mcrdlm1l1_cc_w_1_120_s_3_500=5.02e-12
.param mcrdlm1l1_cf_w_1_120_s_3_500=6.00e-11
.param mcm3m2f_ca_w_0_140_s_0_140=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_140=9.63e-11
.param mcm3m2f_cf_w_0_140_s_0_140=6.58e-12
.param mcm3m2f_ca_w_0_140_s_0_175=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_175=9.45e-11
.param mcm3m2f_cf_w_0_140_s_0_175=8.13e-12
.param mcm3m2f_ca_w_0_140_s_0_210=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_210=8.87e-11
.param mcm3m2f_cf_w_0_140_s_0_210=9.67e-12
.param mcm3m2f_ca_w_0_140_s_0_280=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_280=7.64e-11
.param mcm3m2f_cf_w_0_140_s_0_280=1.26e-11
.param mcm3m2f_ca_w_0_140_s_0_350=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_350=6.46e-11
.param mcm3m2f_cf_w_0_140_s_0_350=1.54e-11
.param mcm3m2f_ca_w_0_140_s_0_420=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_420=5.44e-11
.param mcm3m2f_cf_w_0_140_s_0_420=1.82e-11
.param mcm3m2f_ca_w_0_140_s_0_560=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_560=4.04e-11
.param mcm3m2f_cf_w_0_140_s_0_560=2.31e-11
.param mcm3m2f_ca_w_0_140_s_0_840=9.98e-05
.param mcm3m2f_cc_w_0_140_s_0_840=2.47e-11
.param mcm3m2f_cf_w_0_140_s_0_840=3.11e-11
.param mcm3m2f_ca_w_0_140_s_1_540=9.98e-05
.param mcm3m2f_cc_w_0_140_s_1_540=8.98e-12
.param mcm3m2f_cf_w_0_140_s_1_540=4.26e-11
.param mcm3m2f_ca_w_0_140_s_3_500=9.98e-05
.param mcm3m2f_cc_w_0_140_s_3_500=8.85e-13
.param mcm3m2f_cf_w_0_140_s_3_500=5.01e-11
.param mcm3m2f_ca_w_1_120_s_0_140=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_140=1.08e-10
.param mcm3m2f_cf_w_1_120_s_0_140=6.61e-12
.param mcm3m2f_ca_w_1_120_s_0_175=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_175=1.06e-10
.param mcm3m2f_cf_w_1_120_s_0_175=8.17e-12
.param mcm3m2f_ca_w_1_120_s_0_210=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_210=9.88e-11
.param mcm3m2f_cf_w_1_120_s_0_210=9.69e-12
.param mcm3m2f_ca_w_1_120_s_0_280=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_280=8.46e-11
.param mcm3m2f_cf_w_1_120_s_0_280=1.27e-11
.param mcm3m2f_ca_w_1_120_s_0_350=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_350=7.19e-11
.param mcm3m2f_cf_w_1_120_s_0_350=1.55e-11
.param mcm3m2f_ca_w_1_120_s_0_420=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_420=6.08e-11
.param mcm3m2f_cf_w_1_120_s_0_420=1.82e-11
.param mcm3m2f_ca_w_1_120_s_0_560=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_560=4.53e-11
.param mcm3m2f_cf_w_1_120_s_0_560=2.32e-11
.param mcm3m2f_ca_w_1_120_s_0_840=9.98e-05
.param mcm3m2f_cc_w_1_120_s_0_840=2.81e-11
.param mcm3m2f_cf_w_1_120_s_0_840=3.14e-11
.param mcm3m2f_ca_w_1_120_s_1_540=9.98e-05
.param mcm3m2f_cc_w_1_120_s_1_540=1.07e-11
.param mcm3m2f_cf_w_1_120_s_1_540=4.37e-11
.param mcm3m2f_ca_w_1_120_s_3_500=9.98e-05
.param mcm3m2f_cc_w_1_120_s_3_500=1.09e-12
.param mcm3m2f_cf_w_1_120_s_3_500=5.26e-11
.param mcm3m2d_ca_w_0_140_s_0_140=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_140=9.60e-11
.param mcm3m2d_cf_w_0_140_s_0_140=6.81e-12
.param mcm3m2d_ca_w_0_140_s_0_175=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_175=9.41e-11
.param mcm3m2d_cf_w_0_140_s_0_175=8.42e-12
.param mcm3m2d_ca_w_0_140_s_0_210=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_210=8.84e-11
.param mcm3m2d_cf_w_0_140_s_0_210=1.00e-11
.param mcm3m2d_ca_w_0_140_s_0_280=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_280=7.58e-11
.param mcm3m2d_cf_w_0_140_s_0_280=1.30e-11
.param mcm3m2d_ca_w_0_140_s_0_350=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_350=6.40e-11
.param mcm3m2d_cf_w_0_140_s_0_350=1.60e-11
.param mcm3m2d_ca_w_0_140_s_0_420=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_420=5.36e-11
.param mcm3m2d_cf_w_0_140_s_0_420=1.89e-11
.param mcm3m2d_ca_w_0_140_s_0_560=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_560=3.96e-11
.param mcm3m2d_cf_w_0_140_s_0_560=2.39e-11
.param mcm3m2d_ca_w_0_140_s_0_840=1.03e-04
.param mcm3m2d_cc_w_0_140_s_0_840=2.37e-11
.param mcm3m2d_cf_w_0_140_s_0_840=3.21e-11
.param mcm3m2d_ca_w_0_140_s_1_540=1.03e-04
.param mcm3m2d_cc_w_0_140_s_1_540=8.11e-12
.param mcm3m2d_cf_w_0_140_s_1_540=4.38e-11
.param mcm3m2d_ca_w_0_140_s_3_500=1.03e-04
.param mcm3m2d_cc_w_0_140_s_3_500=6.60e-13
.param mcm3m2d_cf_w_0_140_s_3_500=5.08e-11
.param mcm3m2d_ca_w_1_120_s_0_140=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_140=1.07e-10
.param mcm3m2d_cf_w_1_120_s_0_140=6.85e-12
.param mcm3m2d_ca_w_1_120_s_0_175=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_175=1.05e-10
.param mcm3m2d_cf_w_1_120_s_0_175=8.48e-12
.param mcm3m2d_ca_w_1_120_s_0_210=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_210=9.73e-11
.param mcm3m2d_cf_w_1_120_s_0_210=1.00e-11
.param mcm3m2d_ca_w_1_120_s_0_280=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_280=8.32e-11
.param mcm3m2d_cf_w_1_120_s_0_280=1.31e-11
.param mcm3m2d_ca_w_1_120_s_0_350=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_350=7.03e-11
.param mcm3m2d_cf_w_1_120_s_0_350=1.61e-11
.param mcm3m2d_ca_w_1_120_s_0_420=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_420=5.93e-11
.param mcm3m2d_cf_w_1_120_s_0_420=1.89e-11
.param mcm3m2d_ca_w_1_120_s_0_560=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_560=4.37e-11
.param mcm3m2d_cf_w_1_120_s_0_560=2.41e-11
.param mcm3m2d_ca_w_1_120_s_0_840=1.03e-04
.param mcm3m2d_cc_w_1_120_s_0_840=2.66e-11
.param mcm3m2d_cf_w_1_120_s_0_840=3.25e-11
.param mcm3m2d_ca_w_1_120_s_1_540=1.03e-04
.param mcm3m2d_cc_w_1_120_s_1_540=9.39e-12
.param mcm3m2d_cf_w_1_120_s_1_540=4.48e-11
.param mcm3m2d_ca_w_1_120_s_3_500=1.03e-04
.param mcm3m2d_cc_w_1_120_s_3_500=7.50e-13
.param mcm3m2d_cf_w_1_120_s_3_500=5.30e-11
.param mcm3m2p1_ca_w_0_140_s_0_140=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_140=9.70e-11
.param mcm3m2p1_cf_w_0_140_s_0_140=7.08e-12
.param mcm3m2p1_ca_w_0_140_s_0_175=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_175=9.36e-11
.param mcm3m2p1_cf_w_0_140_s_0_175=8.76e-12
.param mcm3m2p1_ca_w_0_140_s_0_210=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_210=8.75e-11
.param mcm3m2p1_cf_w_0_140_s_0_210=1.04e-11
.param mcm3m2p1_ca_w_0_140_s_0_280=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_280=7.52e-11
.param mcm3m2p1_cf_w_0_140_s_0_280=1.36e-11
.param mcm3m2p1_ca_w_0_140_s_0_350=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_350=6.30e-11
.param mcm3m2p1_cf_w_0_140_s_0_350=1.67e-11
.param mcm3m2p1_ca_w_0_140_s_0_420=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_420=5.27e-11
.param mcm3m2p1_cf_w_0_140_s_0_420=1.96e-11
.param mcm3m2p1_ca_w_0_140_s_0_560=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_560=3.85e-11
.param mcm3m2p1_cf_w_0_140_s_0_560=2.48e-11
.param mcm3m2p1_ca_w_0_140_s_0_840=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_0_840=2.27e-11
.param mcm3m2p1_cf_w_0_140_s_0_840=3.33e-11
.param mcm3m2p1_ca_w_0_140_s_1_540=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_1_540=7.25e-12
.param mcm3m2p1_cf_w_0_140_s_1_540=4.51e-11
.param mcm3m2p1_ca_w_0_140_s_3_500=1.07e-04
.param mcm3m2p1_cc_w_0_140_s_3_500=4.75e-13
.param mcm3m2p1_cf_w_0_140_s_3_500=5.16e-11
.param mcm3m2p1_ca_w_1_120_s_0_140=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_140=1.06e-10
.param mcm3m2p1_cf_w_1_120_s_0_140=7.13e-12
.param mcm3m2p1_ca_w_1_120_s_0_175=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_175=1.03e-10
.param mcm3m2p1_cf_w_1_120_s_0_175=8.82e-12
.param mcm3m2p1_ca_w_1_120_s_0_210=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_210=9.58e-11
.param mcm3m2p1_cf_w_1_120_s_0_210=1.05e-11
.param mcm3m2p1_ca_w_1_120_s_0_280=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_280=8.16e-11
.param mcm3m2p1_cf_w_1_120_s_0_280=1.37e-11
.param mcm3m2p1_ca_w_1_120_s_0_350=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_350=6.87e-11
.param mcm3m2p1_cf_w_1_120_s_0_350=1.68e-11
.param mcm3m2p1_ca_w_1_120_s_0_420=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_420=5.77e-11
.param mcm3m2p1_cf_w_1_120_s_0_420=1.97e-11
.param mcm3m2p1_ca_w_1_120_s_0_560=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_560=4.20e-11
.param mcm3m2p1_cf_w_1_120_s_0_560=2.51e-11
.param mcm3m2p1_ca_w_1_120_s_0_840=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_0_840=2.49e-11
.param mcm3m2p1_cf_w_1_120_s_0_840=3.37e-11
.param mcm3m2p1_ca_w_1_120_s_1_540=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_1_540=8.16e-12
.param mcm3m2p1_cf_w_1_120_s_1_540=4.62e-11
.param mcm3m2p1_ca_w_1_120_s_3_500=1.07e-04
.param mcm3m2p1_cc_w_1_120_s_3_500=5.15e-13
.param mcm3m2p1_cf_w_1_120_s_3_500=5.35e-11
.param mcm3m2l1_ca_w_0_140_s_0_140=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_140=9.45e-11
.param mcm3m2l1_cf_w_0_140_s_0_140=7.89e-12
.param mcm3m2l1_ca_w_0_140_s_0_175=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_175=9.21e-11
.param mcm3m2l1_cf_w_0_140_s_0_175=9.79e-12
.param mcm3m2l1_ca_w_0_140_s_0_210=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_210=8.62e-11
.param mcm3m2l1_cf_w_0_140_s_0_210=1.16e-11
.param mcm3m2l1_ca_w_0_140_s_0_280=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_280=7.32e-11
.param mcm3m2l1_cf_w_0_140_s_0_280=1.52e-11
.param mcm3m2l1_ca_w_0_140_s_0_350=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_350=6.08e-11
.param mcm3m2l1_cf_w_0_140_s_0_350=1.87e-11
.param mcm3m2l1_ca_w_0_140_s_0_420=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_420=5.06e-11
.param mcm3m2l1_cf_w_0_140_s_0_420=2.21e-11
.param mcm3m2l1_ca_w_0_140_s_0_560=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_560=3.58e-11
.param mcm3m2l1_cf_w_0_140_s_0_560=2.78e-11
.param mcm3m2l1_ca_w_0_140_s_0_840=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_0_840=1.98e-11
.param mcm3m2l1_cf_w_0_140_s_0_840=3.71e-11
.param mcm3m2l1_ca_w_0_140_s_1_540=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_1_540=5.20e-12
.param mcm3m2l1_cf_w_0_140_s_1_540=4.89e-11
.param mcm3m2l1_ca_w_0_140_s_3_500=1.19e-04
.param mcm3m2l1_cc_w_0_140_s_3_500=2.10e-13
.param mcm3m2l1_cf_w_0_140_s_3_500=5.38e-11
.param mcm3m2l1_ca_w_1_120_s_0_140=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_140=1.02e-10
.param mcm3m2l1_cf_w_1_120_s_0_140=7.93e-12
.param mcm3m2l1_ca_w_1_120_s_0_175=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_175=9.84e-11
.param mcm3m2l1_cf_w_1_120_s_0_175=9.84e-12
.param mcm3m2l1_ca_w_1_120_s_0_210=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_210=9.19e-11
.param mcm3m2l1_cf_w_1_120_s_0_210=1.17e-11
.param mcm3m2l1_ca_w_1_120_s_0_280=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_280=7.72e-11
.param mcm3m2l1_cf_w_1_120_s_0_280=1.53e-11
.param mcm3m2l1_ca_w_1_120_s_0_350=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_350=6.42e-11
.param mcm3m2l1_cf_w_1_120_s_0_350=1.88e-11
.param mcm3m2l1_ca_w_1_120_s_0_420=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_420=5.32e-11
.param mcm3m2l1_cf_w_1_120_s_0_420=2.21e-11
.param mcm3m2l1_ca_w_1_120_s_0_560=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_560=3.79e-11
.param mcm3m2l1_cf_w_1_120_s_0_560=2.81e-11
.param mcm3m2l1_ca_w_1_120_s_0_840=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_0_840=2.09e-11
.param mcm3m2l1_cf_w_1_120_s_0_840=3.76e-11
.param mcm3m2l1_ca_w_1_120_s_1_540=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_1_540=5.55e-12
.param mcm3m2l1_cf_w_1_120_s_1_540=4.96e-11
.param mcm3m2l1_ca_w_1_120_s_3_500=1.19e-04
.param mcm3m2l1_cc_w_1_120_s_3_500=2.35e-13
.param mcm3m2l1_cf_w_1_120_s_3_500=5.51e-11
.param mcm3m2m1_ca_w_0_140_s_0_140=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_140=8.61e-11
.param mcm3m2m1_cf_w_0_140_s_0_140=1.36e-11
.param mcm3m2m1_ca_w_0_140_s_0_175=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_175=8.31e-11
.param mcm3m2m1_cf_w_0_140_s_0_175=1.70e-11
.param mcm3m2m1_ca_w_0_140_s_0_210=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_210=7.67e-11
.param mcm3m2m1_cf_w_0_140_s_0_210=2.04e-11
.param mcm3m2m1_ca_w_0_140_s_0_280=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_280=6.27e-11
.param mcm3m2m1_cf_w_0_140_s_0_280=2.67e-11
.param mcm3m2m1_ca_w_0_140_s_0_350=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_350=5.02e-11
.param mcm3m2m1_cf_w_0_140_s_0_350=3.24e-11
.param mcm3m2m1_ca_w_0_140_s_0_420=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_420=3.93e-11
.param mcm3m2m1_cf_w_0_140_s_0_420=3.78e-11
.param mcm3m2m1_ca_w_0_140_s_0_560=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_560=2.50e-11
.param mcm3m2m1_cf_w_0_140_s_0_560=4.64e-11
.param mcm3m2m1_ca_w_0_140_s_0_840=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_0_840=1.07e-11
.param mcm3m2m1_cf_w_0_140_s_0_840=5.79e-11
.param mcm3m2m1_ca_w_0_140_s_1_540=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_1_540=1.40e-12
.param mcm3m2m1_cf_w_0_140_s_1_540=6.72e-11
.param mcm3m2m1_ca_w_0_140_s_3_500=2.10e-04
.param mcm3m2m1_cc_w_0_140_s_3_500=3.00e-14
.param mcm3m2m1_cf_w_0_140_s_3_500=6.92e-11
.param mcm3m2m1_ca_w_1_120_s_0_140=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_140=8.88e-11
.param mcm3m2m1_cf_w_1_120_s_0_140=1.36e-11
.param mcm3m2m1_ca_w_1_120_s_0_175=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_175=8.57e-11
.param mcm3m2m1_cf_w_1_120_s_0_175=1.71e-11
.param mcm3m2m1_ca_w_1_120_s_0_210=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_210=7.85e-11
.param mcm3m2m1_cf_w_1_120_s_0_210=2.04e-11
.param mcm3m2m1_ca_w_1_120_s_0_280=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_280=6.38e-11
.param mcm3m2m1_cf_w_1_120_s_0_280=2.67e-11
.param mcm3m2m1_ca_w_1_120_s_0_350=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_350=5.11e-11
.param mcm3m2m1_cf_w_1_120_s_0_350=3.26e-11
.param mcm3m2m1_ca_w_1_120_s_0_420=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_420=4.03e-11
.param mcm3m2m1_cf_w_1_120_s_0_420=3.78e-11
.param mcm3m2m1_ca_w_1_120_s_0_560=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_560=2.57e-11
.param mcm3m2m1_cf_w_1_120_s_0_560=4.67e-11
.param mcm3m2m1_ca_w_1_120_s_0_840=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_0_840=1.09e-11
.param mcm3m2m1_cf_w_1_120_s_0_840=5.84e-11
.param mcm3m2m1_ca_w_1_120_s_1_540=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_1_540=1.40e-12
.param mcm3m2m1_cf_w_1_120_s_1_540=6.78e-11
.param mcm3m2m1_ca_w_1_120_s_3_500=2.10e-04
.param mcm3m2m1_cc_w_1_120_s_3_500=5.00e-14
.param mcm3m2m1_cf_w_1_120_s_3_500=6.98e-11
.param mcm4m2f_ca_w_0_140_s_0_140=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_140=1.04e-10
.param mcm4m2f_cf_w_0_140_s_0_140=2.66e-12
.param mcm4m2f_ca_w_0_140_s_0_175=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_175=1.02e-10
.param mcm4m2f_cf_w_0_140_s_0_175=3.31e-12
.param mcm4m2f_ca_w_0_140_s_0_210=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_210=9.64e-11
.param mcm4m2f_cf_w_0_140_s_0_210=3.98e-12
.param mcm4m2f_ca_w_0_140_s_0_280=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_280=8.50e-11
.param mcm4m2f_cf_w_0_140_s_0_280=5.28e-12
.param mcm4m2f_ca_w_0_140_s_0_350=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_350=7.37e-11
.param mcm4m2f_cf_w_0_140_s_0_350=6.53e-12
.param mcm4m2f_ca_w_0_140_s_0_420=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_420=6.38e-11
.param mcm4m2f_cf_w_0_140_s_0_420=7.86e-12
.param mcm4m2f_ca_w_0_140_s_0_560=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_560=5.04e-11
.param mcm4m2f_cf_w_0_140_s_0_560=1.03e-11
.param mcm4m2f_ca_w_0_140_s_0_840=3.84e-05
.param mcm4m2f_cc_w_0_140_s_0_840=3.52e-11
.param mcm4m2f_cf_w_0_140_s_0_840=1.47e-11
.param mcm4m2f_ca_w_0_140_s_1_540=3.84e-05
.param mcm4m2f_cc_w_0_140_s_1_540=1.76e-11
.param mcm4m2f_cf_w_0_140_s_1_540=2.35e-11
.param mcm4m2f_ca_w_0_140_s_3_500=3.84e-05
.param mcm4m2f_cc_w_0_140_s_3_500=3.53e-12
.param mcm4m2f_cf_w_0_140_s_3_500=3.44e-11
.param mcm4m2f_ca_w_1_120_s_0_140=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_140=1.23e-10
.param mcm4m2f_cf_w_1_120_s_0_140=2.69e-12
.param mcm4m2f_ca_w_1_120_s_0_175=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_175=1.20e-10
.param mcm4m2f_cf_w_1_120_s_0_175=3.34e-12
.param mcm4m2f_ca_w_1_120_s_0_210=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_210=1.13e-10
.param mcm4m2f_cf_w_1_120_s_0_210=4.00e-12
.param mcm4m2f_ca_w_1_120_s_0_280=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_280=9.86e-11
.param mcm4m2f_cf_w_1_120_s_0_280=5.30e-12
.param mcm4m2f_ca_w_1_120_s_0_350=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_350=8.59e-11
.param mcm4m2f_cf_w_1_120_s_0_350=6.58e-12
.param mcm4m2f_ca_w_1_120_s_0_420=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_420=7.50e-11
.param mcm4m2f_cf_w_1_120_s_0_420=7.85e-12
.param mcm4m2f_ca_w_1_120_s_0_560=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_560=5.92e-11
.param mcm4m2f_cf_w_1_120_s_0_560=1.03e-11
.param mcm4m2f_ca_w_1_120_s_0_840=3.84e-05
.param mcm4m2f_cc_w_1_120_s_0_840=4.13e-11
.param mcm4m2f_cf_w_1_120_s_0_840=1.49e-11
.param mcm4m2f_ca_w_1_120_s_1_540=3.84e-05
.param mcm4m2f_cc_w_1_120_s_1_540=2.09e-11
.param mcm4m2f_cf_w_1_120_s_1_540=2.42e-11
.param mcm4m2f_ca_w_1_120_s_3_500=3.84e-05
.param mcm4m2f_cc_w_1_120_s_3_500=4.30e-12
.param mcm4m2f_cf_w_1_120_s_3_500=3.66e-11
.param mcm4m2d_ca_w_0_140_s_0_140=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_140=1.03e-10
.param mcm4m2d_cf_w_0_140_s_0_140=2.89e-12
.param mcm4m2d_ca_w_0_140_s_0_175=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_175=1.01e-10
.param mcm4m2d_cf_w_0_140_s_0_175=3.60e-12
.param mcm4m2d_ca_w_0_140_s_0_210=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_210=9.60e-11
.param mcm4m2d_cf_w_0_140_s_0_210=4.32e-12
.param mcm4m2d_ca_w_0_140_s_0_280=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_280=8.45e-11
.param mcm4m2d_cf_w_0_140_s_0_280=5.73e-12
.param mcm4m2d_ca_w_0_140_s_0_350=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_350=7.30e-11
.param mcm4m2d_cf_w_0_140_s_0_350=7.10e-12
.param mcm4m2d_ca_w_0_140_s_0_420=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_420=6.31e-11
.param mcm4m2d_cf_w_0_140_s_0_420=8.52e-12
.param mcm4m2d_ca_w_0_140_s_0_560=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_560=4.95e-11
.param mcm4m2d_cf_w_0_140_s_0_560=1.11e-11
.param mcm4m2d_ca_w_0_140_s_0_840=4.17e-05
.param mcm4m2d_cc_w_0_140_s_0_840=3.42e-11
.param mcm4m2d_cf_w_0_140_s_0_840=1.59e-11
.param mcm4m2d_ca_w_0_140_s_1_540=4.17e-05
.param mcm4m2d_cc_w_0_140_s_1_540=1.64e-11
.param mcm4m2d_cf_w_0_140_s_1_540=2.51e-11
.param mcm4m2d_ca_w_0_140_s_3_500=4.17e-05
.param mcm4m2d_cc_w_0_140_s_3_500=2.93e-12
.param mcm4m2d_cf_w_0_140_s_3_500=3.60e-11
.param mcm4m2d_ca_w_1_120_s_0_140=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_140=1.22e-10
.param mcm4m2d_cf_w_1_120_s_0_140=2.92e-12
.param mcm4m2d_ca_w_1_120_s_0_175=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_175=1.18e-10
.param mcm4m2d_cf_w_1_120_s_0_175=3.64e-12
.param mcm4m2d_ca_w_1_120_s_0_210=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_210=1.11e-10
.param mcm4m2d_cf_w_1_120_s_0_210=4.35e-12
.param mcm4m2d_ca_w_1_120_s_0_280=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_280=9.72e-11
.param mcm4m2d_cf_w_1_120_s_0_280=5.76e-12
.param mcm4m2d_ca_w_1_120_s_0_350=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_350=8.44e-11
.param mcm4m2d_cf_w_1_120_s_0_350=7.16e-12
.param mcm4m2d_ca_w_1_120_s_0_420=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_420=7.34e-11
.param mcm4m2d_cf_w_1_120_s_0_420=8.53e-12
.param mcm4m2d_ca_w_1_120_s_0_560=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_560=5.76e-11
.param mcm4m2d_cf_w_1_120_s_0_560=1.12e-11
.param mcm4m2d_ca_w_1_120_s_0_840=4.17e-05
.param mcm4m2d_cc_w_1_120_s_0_840=3.96e-11
.param mcm4m2d_cf_w_1_120_s_0_840=1.61e-11
.param mcm4m2d_ca_w_1_120_s_1_540=4.17e-05
.param mcm4m2d_cc_w_1_120_s_1_540=1.93e-11
.param mcm4m2d_cf_w_1_120_s_1_540=2.58e-11
.param mcm4m2d_ca_w_1_120_s_3_500=4.17e-05
.param mcm4m2d_cc_w_1_120_s_3_500=3.51e-12
.param mcm4m2d_cf_w_1_120_s_3_500=3.81e-11
.param mcm4m2p1_ca_w_0_140_s_0_140=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_140=1.03e-10
.param mcm4m2p1_cf_w_0_140_s_0_140=3.16e-12
.param mcm4m2p1_ca_w_0_140_s_0_175=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_175=1.01e-10
.param mcm4m2p1_cf_w_0_140_s_0_175=3.94e-12
.param mcm4m2p1_ca_w_0_140_s_0_210=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_210=9.50e-11
.param mcm4m2p1_cf_w_0_140_s_0_210=4.73e-12
.param mcm4m2p1_ca_w_0_140_s_0_280=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_280=8.37e-11
.param mcm4m2p1_cf_w_0_140_s_0_280=6.26e-12
.param mcm4m2p1_ca_w_0_140_s_0_350=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_350=7.23e-11
.param mcm4m2p1_cf_w_0_140_s_0_350=7.76e-12
.param mcm4m2p1_ca_w_0_140_s_0_420=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_420=6.22e-11
.param mcm4m2p1_cf_w_0_140_s_0_420=9.29e-12
.param mcm4m2p1_ca_w_0_140_s_0_560=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_560=4.88e-11
.param mcm4m2p1_cf_w_0_140_s_0_560=1.21e-11
.param mcm4m2p1_ca_w_0_140_s_0_840=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_0_840=3.29e-11
.param mcm4m2p1_cf_w_0_140_s_0_840=1.72e-11
.param mcm4m2p1_ca_w_0_140_s_1_540=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_1_540=1.52e-11
.param mcm4m2p1_cf_w_0_140_s_1_540=2.69e-11
.param mcm4m2p1_ca_w_0_140_s_3_500=4.56e-05
.param mcm4m2p1_cc_w_0_140_s_3_500=2.39e-12
.param mcm4m2p1_cf_w_0_140_s_3_500=3.75e-11
.param mcm4m2p1_ca_w_1_120_s_0_140=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_140=1.20e-10
.param mcm4m2p1_cf_w_1_120_s_0_140=3.23e-12
.param mcm4m2p1_ca_w_1_120_s_0_175=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_175=1.17e-10
.param mcm4m2p1_cf_w_1_120_s_0_175=4.00e-12
.param mcm4m2p1_ca_w_1_120_s_0_210=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_210=1.10e-10
.param mcm4m2p1_cf_w_1_120_s_0_210=4.77e-12
.param mcm4m2p1_ca_w_1_120_s_0_280=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_280=9.55e-11
.param mcm4m2p1_cf_w_1_120_s_0_280=6.31e-12
.param mcm4m2p1_ca_w_1_120_s_0_350=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_350=8.27e-11
.param mcm4m2p1_cf_w_1_120_s_0_350=7.83e-12
.param mcm4m2p1_ca_w_1_120_s_0_420=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_420=7.18e-11
.param mcm4m2p1_cf_w_1_120_s_0_420=9.33e-12
.param mcm4m2p1_ca_w_1_120_s_0_560=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_560=5.60e-11
.param mcm4m2p1_cf_w_1_120_s_0_560=1.22e-11
.param mcm4m2p1_ca_w_1_120_s_0_840=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_0_840=3.79e-11
.param mcm4m2p1_cf_w_1_120_s_0_840=1.75e-11
.param mcm4m2p1_ca_w_1_120_s_1_540=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_1_540=1.78e-11
.param mcm4m2p1_cf_w_1_120_s_1_540=2.78e-11
.param mcm4m2p1_ca_w_1_120_s_3_500=4.56e-05
.param mcm4m2p1_cc_w_1_120_s_3_500=2.83e-12
.param mcm4m2p1_cf_w_1_120_s_3_500=3.97e-11
.param mcm4m2l1_ca_w_0_140_s_0_140=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_140=1.01e-10
.param mcm4m2l1_cf_w_0_140_s_0_140=3.98e-12
.param mcm4m2l1_ca_w_0_140_s_0_175=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_175=9.91e-11
.param mcm4m2l1_cf_w_0_140_s_0_175=4.97e-12
.param mcm4m2l1_ca_w_0_140_s_0_210=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_210=9.33e-11
.param mcm4m2l1_cf_w_0_140_s_0_210=5.97e-12
.param mcm4m2l1_ca_w_0_140_s_0_280=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_280=8.16e-11
.param mcm4m2l1_cf_w_0_140_s_0_280=7.90e-12
.param mcm4m2l1_ca_w_0_140_s_0_350=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_350=6.99e-11
.param mcm4m2l1_cf_w_0_140_s_0_350=9.78e-12
.param mcm4m2l1_ca_w_0_140_s_0_420=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_420=5.99e-11
.param mcm4m2l1_cf_w_0_140_s_0_420=1.17e-11
.param mcm4m2l1_ca_w_0_140_s_0_560=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_560=4.60e-11
.param mcm4m2l1_cf_w_0_140_s_0_560=1.52e-11
.param mcm4m2l1_ca_w_0_140_s_0_840=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_0_840=2.99e-11
.param mcm4m2l1_cf_w_0_140_s_0_840=2.13e-11
.param mcm4m2l1_ca_w_0_140_s_1_540=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_1_540=1.24e-11
.param mcm4m2l1_cf_w_0_140_s_1_540=3.21e-11
.param mcm4m2l1_ca_w_0_140_s_3_500=5.79e-05
.param mcm4m2l1_cc_w_0_140_s_3_500=1.46e-12
.param mcm4m2l1_cf_w_0_140_s_3_500=4.17e-11
.param mcm4m2l1_ca_w_1_120_s_0_140=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_140=1.16e-10
.param mcm4m2l1_cf_w_1_120_s_0_140=4.01e-12
.param mcm4m2l1_ca_w_1_120_s_0_175=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_175=1.13e-10
.param mcm4m2l1_cf_w_1_120_s_0_175=5.01e-12
.param mcm4m2l1_ca_w_1_120_s_0_210=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_210=1.06e-10
.param mcm4m2l1_cf_w_1_120_s_0_210=6.00e-12
.param mcm4m2l1_ca_w_1_120_s_0_280=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_280=9.13e-11
.param mcm4m2l1_cf_w_1_120_s_0_280=7.94e-12
.param mcm4m2l1_ca_w_1_120_s_0_350=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_350=7.86e-11
.param mcm4m2l1_cf_w_1_120_s_0_350=9.87e-12
.param mcm4m2l1_ca_w_1_120_s_0_420=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_420=6.73e-11
.param mcm4m2l1_cf_w_1_120_s_0_420=1.17e-11
.param mcm4m2l1_ca_w_1_120_s_0_560=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_560=5.17e-11
.param mcm4m2l1_cf_w_1_120_s_0_560=1.52e-11
.param mcm4m2l1_ca_w_1_120_s_0_840=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_0_840=3.38e-11
.param mcm4m2l1_cf_w_1_120_s_0_840=2.16e-11
.param mcm4m2l1_ca_w_1_120_s_1_540=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_1_540=1.44e-11
.param mcm4m2l1_cf_w_1_120_s_1_540=3.30e-11
.param mcm4m2l1_ca_w_1_120_s_3_500=5.79e-05
.param mcm4m2l1_cc_w_1_120_s_3_500=1.71e-12
.param mcm4m2l1_cf_w_1_120_s_3_500=4.38e-11
.param mcm4m2m1_ca_w_0_140_s_0_140=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_140=9.29e-11
.param mcm4m2m1_cf_w_0_140_s_0_140=9.69e-12
.param mcm4m2m1_ca_w_0_140_s_0_175=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_175=9.05e-11
.param mcm4m2m1_cf_w_0_140_s_0_175=1.22e-11
.param mcm4m2m1_ca_w_0_140_s_0_210=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_210=8.43e-11
.param mcm4m2m1_cf_w_0_140_s_0_210=1.47e-11
.param mcm4m2m1_ca_w_0_140_s_0_280=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_280=7.12e-11
.param mcm4m2m1_cf_w_0_140_s_0_280=1.93e-11
.param mcm4m2m1_ca_w_0_140_s_0_350=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_350=5.89e-11
.param mcm4m2m1_cf_w_0_140_s_0_350=2.36e-11
.param mcm4m2m1_ca_w_0_140_s_0_420=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_420=4.87e-11
.param mcm4m2m1_cf_w_0_140_s_0_420=2.76e-11
.param mcm4m2m1_ca_w_0_140_s_0_560=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_560=3.47e-11
.param mcm4m2m1_cf_w_0_140_s_0_560=3.43e-11
.param mcm4m2m1_ca_w_0_140_s_0_840=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_0_840=1.95e-11
.param mcm4m2m1_cf_w_0_140_s_0_840=4.42e-11
.param mcm4m2m1_ca_w_0_140_s_1_540=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_1_540=5.90e-12
.param mcm4m2m1_cf_w_0_140_s_1_540=5.59e-11
.param mcm4m2m1_ca_w_0_140_s_3_500=1.49e-04
.param mcm4m2m1_cc_w_0_140_s_3_500=3.95e-13
.param mcm4m2m1_cf_w_0_140_s_3_500=6.18e-11
.param mcm4m2m1_ca_w_1_120_s_0_140=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_140=1.02e-10
.param mcm4m2m1_cf_w_1_120_s_0_140=9.67e-12
.param mcm4m2m1_ca_w_1_120_s_0_175=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_175=9.96e-11
.param mcm4m2m1_cf_w_1_120_s_0_175=1.22e-11
.param mcm4m2m1_ca_w_1_120_s_0_210=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_210=9.26e-11
.param mcm4m2m1_cf_w_1_120_s_0_210=1.47e-11
.param mcm4m2m1_ca_w_1_120_s_0_280=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_280=7.82e-11
.param mcm4m2m1_cf_w_1_120_s_0_280=1.93e-11
.param mcm4m2m1_ca_w_1_120_s_0_350=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_350=6.51e-11
.param mcm4m2m1_cf_w_1_120_s_0_350=2.36e-11
.param mcm4m2m1_ca_w_1_120_s_0_420=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_420=5.43e-11
.param mcm4m2m1_cf_w_1_120_s_0_420=2.76e-11
.param mcm4m2m1_ca_w_1_120_s_0_560=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_560=3.91e-11
.param mcm4m2m1_cf_w_1_120_s_0_560=3.44e-11
.param mcm4m2m1_ca_w_1_120_s_0_840=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_0_840=2.27e-11
.param mcm4m2m1_cf_w_1_120_s_0_840=4.46e-11
.param mcm4m2m1_ca_w_1_120_s_1_540=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_1_540=7.30e-12
.param mcm4m2m1_cf_w_1_120_s_1_540=5.73e-11
.param mcm4m2m1_ca_w_1_120_s_3_500=1.49e-04
.param mcm4m2m1_cc_w_1_120_s_3_500=5.30e-13
.param mcm4m2m1_cf_w_1_120_s_3_500=6.42e-11
.param mcm5m2f_ca_w_0_140_s_0_140=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_140=1.05e-10
.param mcm5m2f_cf_w_0_140_s_0_140=2.02e-12
.param mcm5m2f_ca_w_0_140_s_0_175=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_175=1.03e-10
.param mcm5m2f_cf_w_0_140_s_0_175=2.52e-12
.param mcm5m2f_ca_w_0_140_s_0_210=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_210=9.74e-11
.param mcm5m2f_cf_w_0_140_s_0_210=3.03e-12
.param mcm5m2f_ca_w_0_140_s_0_280=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_280=8.66e-11
.param mcm5m2f_cf_w_0_140_s_0_280=4.03e-12
.param mcm5m2f_ca_w_0_140_s_0_350=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_350=7.55e-11
.param mcm5m2f_cf_w_0_140_s_0_350=5.00e-12
.param mcm5m2f_ca_w_0_140_s_0_420=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_420=6.59e-11
.param mcm5m2f_cf_w_0_140_s_0_420=6.02e-12
.param mcm5m2f_ca_w_0_140_s_0_560=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_560=5.27e-11
.param mcm5m2f_cf_w_0_140_s_0_560=7.88e-12
.param mcm5m2f_ca_w_0_140_s_0_840=2.91e-05
.param mcm5m2f_cc_w_0_140_s_0_840=3.83e-11
.param mcm5m2f_cf_w_0_140_s_0_840=1.14e-11
.param mcm5m2f_ca_w_0_140_s_1_540=2.91e-05
.param mcm5m2f_cc_w_0_140_s_1_540=2.12e-11
.param mcm5m2f_cf_w_0_140_s_1_540=1.88e-11
.param mcm5m2f_ca_w_0_140_s_3_500=2.91e-05
.param mcm5m2f_cc_w_0_140_s_3_500=5.84e-12
.param mcm5m2f_cf_w_0_140_s_3_500=2.97e-11
.param mcm5m2f_ca_w_1_120_s_0_140=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_140=1.27e-10
.param mcm5m2f_cf_w_1_120_s_0_140=2.04e-12
.param mcm5m2f_ca_w_1_120_s_0_175=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_175=1.24e-10
.param mcm5m2f_cf_w_1_120_s_0_175=2.55e-12
.param mcm5m2f_ca_w_1_120_s_0_210=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_210=1.17e-10
.param mcm5m2f_cf_w_1_120_s_0_210=3.05e-12
.param mcm5m2f_ca_w_1_120_s_0_280=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_280=1.03e-10
.param mcm5m2f_cf_w_1_120_s_0_280=4.05e-12
.param mcm5m2f_ca_w_1_120_s_0_350=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_350=9.06e-11
.param mcm5m2f_cf_w_1_120_s_0_350=5.03e-12
.param mcm5m2f_ca_w_1_120_s_0_420=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_420=7.97e-11
.param mcm5m2f_cf_w_1_120_s_0_420=6.03e-12
.param mcm5m2f_ca_w_1_120_s_0_560=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_560=6.41e-11
.param mcm5m2f_cf_w_1_120_s_0_560=7.91e-12
.param mcm5m2f_ca_w_1_120_s_0_840=2.91e-05
.param mcm5m2f_cc_w_1_120_s_0_840=4.63e-11
.param mcm5m2f_cf_w_1_120_s_0_840=1.15e-11
.param mcm5m2f_ca_w_1_120_s_1_540=2.91e-05
.param mcm5m2f_cc_w_1_120_s_1_540=2.59e-11
.param mcm5m2f_cf_w_1_120_s_1_540=1.92e-11
.param mcm5m2f_ca_w_1_120_s_3_500=2.91e-05
.param mcm5m2f_cc_w_1_120_s_3_500=7.36e-12
.param mcm5m2f_cf_w_1_120_s_3_500=3.17e-11
.param mcm5m2d_ca_w_0_140_s_0_140=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_140=1.05e-10
.param mcm5m2d_cf_w_0_140_s_0_140=2.25e-12
.param mcm5m2d_ca_w_0_140_s_0_175=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_175=1.02e-10
.param mcm5m2d_cf_w_0_140_s_0_175=2.81e-12
.param mcm5m2d_ca_w_0_140_s_0_210=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_210=9.70e-11
.param mcm5m2d_cf_w_0_140_s_0_210=3.37e-12
.param mcm5m2d_ca_w_0_140_s_0_280=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_280=8.61e-11
.param mcm5m2d_cf_w_0_140_s_0_280=4.48e-12
.param mcm5m2d_ca_w_0_140_s_0_350=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_350=7.48e-11
.param mcm5m2d_cf_w_0_140_s_0_350=5.57e-12
.param mcm5m2d_ca_w_0_140_s_0_420=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_420=6.50e-11
.param mcm5m2d_cf_w_0_140_s_0_420=6.67e-12
.param mcm5m2d_ca_w_0_140_s_0_560=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_560=5.20e-11
.param mcm5m2d_cf_w_0_140_s_0_560=8.75e-12
.param mcm5m2d_ca_w_0_140_s_0_840=3.23e-05
.param mcm5m2d_cc_w_0_140_s_0_840=3.73e-11
.param mcm5m2d_cf_w_0_140_s_0_840=1.26e-11
.param mcm5m2d_ca_w_0_140_s_1_540=3.23e-05
.param mcm5m2d_cc_w_0_140_s_1_540=1.99e-11
.param mcm5m2d_cf_w_0_140_s_1_540=2.05e-11
.param mcm5m2d_ca_w_0_140_s_3_500=3.23e-05
.param mcm5m2d_cc_w_0_140_s_3_500=5.02e-12
.param mcm5m2d_cf_w_0_140_s_3_500=3.15e-11
.param mcm5m2d_ca_w_1_120_s_0_140=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_140=1.26e-10
.param mcm5m2d_cf_w_1_120_s_0_140=2.28e-12
.param mcm5m2d_ca_w_1_120_s_0_175=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_175=1.23e-10
.param mcm5m2d_cf_w_1_120_s_0_175=2.85e-12
.param mcm5m2d_ca_w_1_120_s_0_210=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_210=1.16e-10
.param mcm5m2d_cf_w_1_120_s_0_210=3.40e-12
.param mcm5m2d_ca_w_1_120_s_0_280=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_280=1.02e-10
.param mcm5m2d_cf_w_1_120_s_0_280=4.51e-12
.param mcm5m2d_ca_w_1_120_s_0_350=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_350=8.90e-11
.param mcm5m2d_cf_w_1_120_s_0_350=5.61e-12
.param mcm5m2d_ca_w_1_120_s_0_420=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_420=7.81e-11
.param mcm5m2d_cf_w_1_120_s_0_420=6.69e-12
.param mcm5m2d_ca_w_1_120_s_0_560=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_560=6.25e-11
.param mcm5m2d_cf_w_1_120_s_0_560=8.79e-12
.param mcm5m2d_ca_w_1_120_s_0_840=3.23e-05
.param mcm5m2d_cc_w_1_120_s_0_840=4.46e-11
.param mcm5m2d_cf_w_1_120_s_0_840=1.28e-11
.param mcm5m2d_ca_w_1_120_s_1_540=3.23e-05
.param mcm5m2d_cc_w_1_120_s_1_540=2.43e-11
.param mcm5m2d_cf_w_1_120_s_1_540=2.11e-11
.param mcm5m2d_ca_w_1_120_s_3_500=3.23e-05
.param mcm5m2d_cc_w_1_120_s_3_500=6.40e-12
.param mcm5m2d_cf_w_1_120_s_3_500=3.37e-11
.param mcm5m2p1_ca_w_0_140_s_0_140=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_140=1.04e-10
.param mcm5m2p1_cf_w_0_140_s_0_140=2.52e-12
.param mcm5m2p1_ca_w_0_140_s_0_175=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_175=1.02e-10
.param mcm5m2p1_cf_w_0_140_s_0_175=3.15e-12
.param mcm5m2p1_ca_w_0_140_s_0_210=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_210=9.64e-11
.param mcm5m2p1_cf_w_0_140_s_0_210=3.78e-12
.param mcm5m2p1_ca_w_0_140_s_0_280=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_280=8.54e-11
.param mcm5m2p1_cf_w_0_140_s_0_280=5.02e-12
.param mcm5m2p1_ca_w_0_140_s_0_350=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_350=7.35e-11
.param mcm5m2p1_cf_w_0_140_s_0_350=6.23e-12
.param mcm5m2p1_ca_w_0_140_s_0_420=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_420=6.42e-11
.param mcm5m2p1_cf_w_0_140_s_0_420=7.45e-12
.param mcm5m2p1_ca_w_0_140_s_0_560=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_560=5.11e-11
.param mcm5m2p1_cf_w_0_140_s_0_560=9.75e-12
.param mcm5m2p1_ca_w_0_140_s_0_840=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_0_840=3.60e-11
.param mcm5m2p1_cf_w_0_140_s_0_840=1.40e-11
.param mcm5m2p1_ca_w_0_140_s_1_540=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_1_540=1.87e-11
.param mcm5m2p1_cf_w_0_140_s_1_540=2.25e-11
.param mcm5m2p1_ca_w_0_140_s_3_500=3.62e-05
.param mcm5m2p1_cc_w_0_140_s_3_500=4.31e-12
.param mcm5m2p1_cf_w_0_140_s_3_500=3.34e-11
.param mcm5m2p1_ca_w_1_120_s_0_140=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_140=1.24e-10
.param mcm5m2p1_cf_w_1_120_s_0_140=2.59e-12
.param mcm5m2p1_ca_w_1_120_s_0_175=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_175=1.20e-10
.param mcm5m2p1_cf_w_1_120_s_0_175=3.22e-12
.param mcm5m2p1_ca_w_1_120_s_0_210=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_210=1.14e-10
.param mcm5m2p1_cf_w_1_120_s_0_210=3.85e-12
.param mcm5m2p1_ca_w_1_120_s_0_280=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_280=1.00e-10
.param mcm5m2p1_cf_w_1_120_s_0_280=5.07e-12
.param mcm5m2p1_ca_w_1_120_s_0_350=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_350=8.73e-11
.param mcm5m2p1_cf_w_1_120_s_0_350=6.28e-12
.param mcm5m2p1_ca_w_1_120_s_0_420=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_420=7.65e-11
.param mcm5m2p1_cf_w_1_120_s_0_420=7.49e-12
.param mcm5m2p1_ca_w_1_120_s_0_560=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_560=6.08e-11
.param mcm5m2p1_cf_w_1_120_s_0_560=9.82e-12
.param mcm5m2p1_ca_w_1_120_s_0_840=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_0_840=4.29e-11
.param mcm5m2p1_cf_w_1_120_s_0_840=1.42e-11
.param mcm5m2p1_ca_w_1_120_s_1_540=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_1_540=2.26e-11
.param mcm5m2p1_cf_w_1_120_s_1_540=2.31e-11
.param mcm5m2p1_ca_w_1_120_s_3_500=3.62e-05
.param mcm5m2p1_cc_w_1_120_s_3_500=5.47e-12
.param mcm5m2p1_cf_w_1_120_s_3_500=3.58e-11
.param mcm5m2l1_ca_w_0_140_s_0_140=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_140=1.02e-10
.param mcm5m2l1_cf_w_0_140_s_0_140=3.34e-12
.param mcm5m2l1_ca_w_0_140_s_0_175=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_175=1.00e-10
.param mcm5m2l1_cf_w_0_140_s_0_175=4.18e-12
.param mcm5m2l1_ca_w_0_140_s_0_210=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_210=9.47e-11
.param mcm5m2l1_cf_w_0_140_s_0_210=5.02e-12
.param mcm5m2l1_ca_w_0_140_s_0_280=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_280=8.34e-11
.param mcm5m2l1_cf_w_0_140_s_0_280=6.66e-12
.param mcm5m2l1_ca_w_0_140_s_0_350=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_350=7.14e-11
.param mcm5m2l1_cf_w_0_140_s_0_350=8.25e-12
.param mcm5m2l1_ca_w_0_140_s_0_420=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_420=6.13e-11
.param mcm5m2l1_cf_w_0_140_s_0_420=9.85e-12
.param mcm5m2l1_ca_w_0_140_s_0_560=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_560=4.83e-11
.param mcm5m2l1_cf_w_0_140_s_0_560=1.28e-11
.param mcm5m2l1_ca_w_0_140_s_0_840=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_0_840=3.27e-11
.param mcm5m2l1_cf_w_0_140_s_0_840=1.81e-11
.param mcm5m2l1_ca_w_0_140_s_1_540=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_1_540=1.56e-11
.param mcm5m2l1_cf_w_0_140_s_1_540=2.80e-11
.param mcm5m2l1_ca_w_0_140_s_3_500=4.85e-05
.param mcm5m2l1_cc_w_0_140_s_3_500=2.91e-12
.param mcm5m2l1_cf_w_0_140_s_3_500=3.85e-11
.param mcm5m2l1_ca_w_1_120_s_0_140=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_140=1.20e-10
.param mcm5m2l1_cf_w_1_120_s_0_140=3.37e-12
.param mcm5m2l1_ca_w_1_120_s_0_175=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_175=1.17e-10
.param mcm5m2l1_cf_w_1_120_s_0_175=4.22e-12
.param mcm5m2l1_ca_w_1_120_s_0_210=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_210=1.10e-10
.param mcm5m2l1_cf_w_1_120_s_0_210=5.05e-12
.param mcm5m2l1_ca_w_1_120_s_0_280=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_280=9.58e-11
.param mcm5m2l1_cf_w_1_120_s_0_280=6.69e-12
.param mcm5m2l1_ca_w_1_120_s_0_350=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_350=8.29e-11
.param mcm5m2l1_cf_w_1_120_s_0_350=8.30e-12
.param mcm5m2l1_ca_w_1_120_s_0_420=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_420=7.19e-11
.param mcm5m2l1_cf_w_1_120_s_0_420=9.87e-12
.param mcm5m2l1_ca_w_1_120_s_0_560=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_560=5.65e-11
.param mcm5m2l1_cf_w_1_120_s_0_560=1.29e-11
.param mcm5m2l1_ca_w_1_120_s_0_840=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_0_840=3.88e-11
.param mcm5m2l1_cf_w_1_120_s_0_840=1.83e-11
.param mcm5m2l1_ca_w_1_120_s_1_540=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_1_540=1.90e-11
.param mcm5m2l1_cf_w_1_120_s_1_540=2.87e-11
.param mcm5m2l1_ca_w_1_120_s_3_500=4.85e-05
.param mcm5m2l1_cc_w_1_120_s_3_500=3.81e-12
.param mcm5m2l1_cf_w_1_120_s_3_500=4.09e-11
.param mcm5m2m1_ca_w_0_140_s_0_140=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_140=9.44e-11
.param mcm5m2m1_cf_w_0_140_s_0_140=9.06e-12
.param mcm5m2m1_ca_w_0_140_s_0_175=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_175=9.18e-11
.param mcm5m2m1_cf_w_0_140_s_0_175=1.14e-11
.param mcm5m2m1_ca_w_0_140_s_0_210=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_210=8.57e-11
.param mcm5m2m1_cf_w_0_140_s_0_210=1.37e-11
.param mcm5m2m1_ca_w_0_140_s_0_280=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_280=7.29e-11
.param mcm5m2m1_cf_w_0_140_s_0_280=1.81e-11
.param mcm5m2m1_ca_w_0_140_s_0_350=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_350=6.06e-11
.param mcm5m2m1_cf_w_0_140_s_0_350=2.20e-11
.param mcm5m2m1_ca_w_0_140_s_0_420=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_420=5.08e-11
.param mcm5m2m1_cf_w_0_140_s_0_420=2.58e-11
.param mcm5m2m1_ca_w_0_140_s_0_560=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_560=3.70e-11
.param mcm5m2m1_cf_w_0_140_s_0_560=3.20e-11
.param mcm5m2m1_ca_w_0_140_s_0_840=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_0_840=2.21e-11
.param mcm5m2m1_cf_w_0_140_s_0_840=4.14e-11
.param mcm5m2m1_ca_w_0_140_s_1_540=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_1_540=8.08e-12
.param mcm5m2m1_cf_w_0_140_s_1_540=5.33e-11
.param mcm5m2m1_ca_w_0_140_s_3_500=1.39e-04
.param mcm5m2m1_cc_w_0_140_s_3_500=1.04e-12
.param mcm5m2m1_cf_w_0_140_s_3_500=6.04e-11
.param mcm5m2m1_ca_w_1_120_s_0_140=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_140=1.06e-10
.param mcm5m2m1_cf_w_1_120_s_0_140=9.04e-12
.param mcm5m2m1_ca_w_1_120_s_0_175=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_175=1.03e-10
.param mcm5m2m1_cf_w_1_120_s_0_175=1.15e-11
.param mcm5m2m1_ca_w_1_120_s_0_210=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_210=9.69e-11
.param mcm5m2m1_cf_w_1_120_s_0_210=1.37e-11
.param mcm5m2m1_ca_w_1_120_s_0_280=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_280=8.26e-11
.param mcm5m2m1_cf_w_1_120_s_0_280=1.80e-11
.param mcm5m2m1_ca_w_1_120_s_0_350=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_350=6.94e-11
.param mcm5m2m1_cf_w_1_120_s_0_350=2.20e-11
.param mcm5m2m1_ca_w_1_120_s_0_420=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_420=5.87e-11
.param mcm5m2m1_cf_w_1_120_s_0_420=2.57e-11
.param mcm5m2m1_ca_w_1_120_s_0_560=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_560=4.37e-11
.param mcm5m2m1_cf_w_1_120_s_0_560=3.20e-11
.param mcm5m2m1_ca_w_1_120_s_0_840=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_0_840=2.73e-11
.param mcm5m2m1_cf_w_1_120_s_0_840=4.17e-11
.param mcm5m2m1_ca_w_1_120_s_1_540=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_1_540=1.10e-11
.param mcm5m2m1_cf_w_1_120_s_1_540=5.46e-11
.param mcm5m2m1_ca_w_1_120_s_3_500=1.39e-04
.param mcm5m2m1_cc_w_1_120_s_3_500=1.59e-12
.param mcm5m2m1_cf_w_1_120_s_3_500=6.38e-11
.param mcrdlm2f_ca_w_0_140_s_0_140=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_140=1.06e-10
.param mcrdlm2f_cf_w_0_140_s_0_140=1.44e-12
.param mcrdlm2f_ca_w_0_140_s_0_175=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_175=1.04e-10
.param mcrdlm2f_cf_w_0_140_s_0_175=1.80e-12
.param mcrdlm2f_ca_w_0_140_s_0_210=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_210=9.87e-11
.param mcrdlm2f_cf_w_0_140_s_0_210=2.16e-12
.param mcrdlm2f_ca_w_0_140_s_0_280=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_280=8.79e-11
.param mcrdlm2f_cf_w_0_140_s_0_280=2.88e-12
.param mcrdlm2f_ca_w_0_140_s_0_350=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_350=7.66e-11
.param mcrdlm2f_cf_w_0_140_s_0_350=3.58e-12
.param mcrdlm2f_ca_w_0_140_s_0_420=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_420=6.79e-11
.param mcrdlm2f_cf_w_0_140_s_0_420=4.31e-12
.param mcrdlm2f_ca_w_0_140_s_0_560=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_560=5.51e-11
.param mcrdlm2f_cf_w_0_140_s_0_560=5.64e-12
.param mcrdlm2f_ca_w_0_140_s_0_840=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_0_840=4.14e-11
.param mcrdlm2f_cf_w_0_140_s_0_840=8.21e-12
.param mcrdlm2f_ca_w_0_140_s_1_540=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_1_540=2.56e-11
.param mcrdlm2f_cf_w_0_140_s_1_540=1.39e-11
.param mcrdlm2f_ca_w_0_140_s_3_500=2.06e-05
.param mcrdlm2f_cc_w_0_140_s_3_500=1.02e-11
.param mcrdlm2f_cf_w_0_140_s_3_500=2.38e-11
.param mcrdlm2f_ca_w_1_120_s_0_140=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_140=1.32e-10
.param mcrdlm2f_cf_w_1_120_s_0_140=1.48e-12
.param mcrdlm2f_ca_w_1_120_s_0_175=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_175=1.28e-10
.param mcrdlm2f_cf_w_1_120_s_0_175=1.84e-12
.param mcrdlm2f_ca_w_1_120_s_0_210=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_210=1.22e-10
.param mcrdlm2f_cf_w_1_120_s_0_210=2.20e-12
.param mcrdlm2f_ca_w_1_120_s_0_280=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_280=1.08e-10
.param mcrdlm2f_cf_w_1_120_s_0_280=2.91e-12
.param mcrdlm2f_ca_w_1_120_s_0_350=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_350=9.52e-11
.param mcrdlm2f_cf_w_1_120_s_0_350=3.62e-12
.param mcrdlm2f_ca_w_1_120_s_0_420=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_420=8.46e-11
.param mcrdlm2f_cf_w_1_120_s_0_420=4.32e-12
.param mcrdlm2f_ca_w_1_120_s_0_560=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_560=6.97e-11
.param mcrdlm2f_cf_w_1_120_s_0_560=5.68e-12
.param mcrdlm2f_ca_w_1_120_s_0_840=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_0_840=5.25e-11
.param mcrdlm2f_cf_w_1_120_s_0_840=8.31e-12
.param mcrdlm2f_ca_w_1_120_s_1_540=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_1_540=3.30e-11
.param mcrdlm2f_cf_w_1_120_s_1_540=1.42e-11
.param mcrdlm2f_ca_w_1_120_s_3_500=2.06e-05
.param mcrdlm2f_cc_w_1_120_s_3_500=1.39e-11
.param mcrdlm2f_cf_w_1_120_s_3_500=2.53e-11
.param mcrdlm2d_ca_w_0_140_s_0_140=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_140=1.05e-10
.param mcrdlm2d_cf_w_0_140_s_0_140=1.67e-12
.param mcrdlm2d_ca_w_0_140_s_0_175=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_175=1.04e-10
.param mcrdlm2d_cf_w_0_140_s_0_175=2.08e-12
.param mcrdlm2d_ca_w_0_140_s_0_210=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_210=9.82e-11
.param mcrdlm2d_cf_w_0_140_s_0_210=2.51e-12
.param mcrdlm2d_ca_w_0_140_s_0_280=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_280=8.74e-11
.param mcrdlm2d_cf_w_0_140_s_0_280=3.33e-12
.param mcrdlm2d_ca_w_0_140_s_0_350=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_350=7.60e-11
.param mcrdlm2d_cf_w_0_140_s_0_350=4.14e-12
.param mcrdlm2d_ca_w_0_140_s_0_420=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_420=6.72e-11
.param mcrdlm2d_cf_w_0_140_s_0_420=4.98e-12
.param mcrdlm2d_ca_w_0_140_s_0_560=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_560=5.42e-11
.param mcrdlm2d_cf_w_0_140_s_0_560=6.50e-12
.param mcrdlm2d_ca_w_0_140_s_0_840=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_0_840=4.02e-11
.param mcrdlm2d_cf_w_0_140_s_0_840=9.43e-12
.param mcrdlm2d_ca_w_0_140_s_1_540=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_1_540=2.42e-11
.param mcrdlm2d_cf_w_0_140_s_1_540=1.57e-11
.param mcrdlm2d_ca_w_0_140_s_3_500=2.39e-05
.param mcrdlm2d_cc_w_0_140_s_3_500=9.06e-12
.param mcrdlm2d_cf_w_0_140_s_3_500=2.61e-11
.param mcrdlm2d_ca_w_1_120_s_0_140=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_140=1.30e-10
.param mcrdlm2d_cf_w_1_120_s_0_140=1.71e-12
.param mcrdlm2d_ca_w_1_120_s_0_175=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_175=1.26e-10
.param mcrdlm2d_cf_w_1_120_s_0_175=2.13e-12
.param mcrdlm2d_ca_w_1_120_s_0_210=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_210=1.20e-10
.param mcrdlm2d_cf_w_1_120_s_0_210=2.55e-12
.param mcrdlm2d_ca_w_1_120_s_0_280=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_280=1.06e-10
.param mcrdlm2d_cf_w_1_120_s_0_280=3.37e-12
.param mcrdlm2d_ca_w_1_120_s_0_350=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_350=9.41e-11
.param mcrdlm2d_cf_w_1_120_s_0_350=4.19e-12
.param mcrdlm2d_ca_w_1_120_s_0_420=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_420=8.30e-11
.param mcrdlm2d_cf_w_1_120_s_0_420=4.99e-12
.param mcrdlm2d_ca_w_1_120_s_0_560=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_560=6.81e-11
.param mcrdlm2d_cf_w_1_120_s_0_560=6.56e-12
.param mcrdlm2d_ca_w_1_120_s_0_840=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_0_840=5.07e-11
.param mcrdlm2d_cf_w_1_120_s_0_840=9.53e-12
.param mcrdlm2d_ca_w_1_120_s_1_540=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_1_540=3.12e-11
.param mcrdlm2d_cf_w_1_120_s_1_540=1.61e-11
.param mcrdlm2d_ca_w_1_120_s_3_500=2.39e-05
.param mcrdlm2d_cc_w_1_120_s_3_500=1.26e-11
.param mcrdlm2d_cf_w_1_120_s_3_500=2.78e-11
.param mcrdlm2p1_ca_w_0_140_s_0_140=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_140=1.05e-10
.param mcrdlm2p1_cf_w_0_140_s_0_140=1.94e-12
.param mcrdlm2p1_ca_w_0_140_s_0_175=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_175=1.03e-10
.param mcrdlm2p1_cf_w_0_140_s_0_175=2.42e-12
.param mcrdlm2p1_ca_w_0_140_s_0_210=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_210=9.76e-11
.param mcrdlm2p1_cf_w_0_140_s_0_210=2.91e-12
.param mcrdlm2p1_ca_w_0_140_s_0_280=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_280=8.67e-11
.param mcrdlm2p1_cf_w_0_140_s_0_280=3.86e-12
.param mcrdlm2p1_ca_w_0_140_s_0_350=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_350=7.54e-11
.param mcrdlm2p1_cf_w_0_140_s_0_350=4.79e-12
.param mcrdlm2p1_ca_w_0_140_s_0_420=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_420=6.64e-11
.param mcrdlm2p1_cf_w_0_140_s_0_420=5.76e-12
.param mcrdlm2p1_ca_w_0_140_s_0_560=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_560=5.33e-11
.param mcrdlm2p1_cf_w_0_140_s_0_560=7.53e-12
.param mcrdlm2p1_ca_w_0_140_s_0_840=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_0_840=3.90e-11
.param mcrdlm2p1_cf_w_0_140_s_0_840=1.09e-11
.param mcrdlm2p1_ca_w_0_140_s_1_540=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_1_540=2.28e-11
.param mcrdlm2p1_cf_w_0_140_s_1_540=1.78e-11
.param mcrdlm2p1_ca_w_0_140_s_3_500=2.78e-05
.param mcrdlm2p1_cc_w_0_140_s_3_500=8.01e-12
.param mcrdlm2p1_cf_w_0_140_s_3_500=2.86e-11
.param mcrdlm2p1_ca_w_1_120_s_0_140=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_140=1.29e-10
.param mcrdlm2p1_cf_w_1_120_s_0_140=2.02e-12
.param mcrdlm2p1_ca_w_1_120_s_0_175=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_175=1.25e-10
.param mcrdlm2p1_cf_w_1_120_s_0_175=2.49e-12
.param mcrdlm2p1_ca_w_1_120_s_0_210=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_210=1.19e-10
.param mcrdlm2p1_cf_w_1_120_s_0_210=2.97e-12
.param mcrdlm2p1_ca_w_1_120_s_0_280=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_280=1.05e-10
.param mcrdlm2p1_cf_w_1_120_s_0_280=3.92e-12
.param mcrdlm2p1_ca_w_1_120_s_0_350=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_350=9.25e-11
.param mcrdlm2p1_cf_w_1_120_s_0_350=4.87e-12
.param mcrdlm2p1_ca_w_1_120_s_0_420=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_420=8.15e-11
.param mcrdlm2p1_cf_w_1_120_s_0_420=5.79e-12
.param mcrdlm2p1_ca_w_1_120_s_0_560=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_560=6.62e-11
.param mcrdlm2p1_cf_w_1_120_s_0_560=7.60e-12
.param mcrdlm2p1_ca_w_1_120_s_0_840=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_0_840=4.91e-11
.param mcrdlm2p1_cf_w_1_120_s_0_840=1.10e-11
.param mcrdlm2p1_ca_w_1_120_s_1_540=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_1_540=2.95e-11
.param mcrdlm2p1_cf_w_1_120_s_1_540=1.82e-11
.param mcrdlm2p1_ca_w_1_120_s_3_500=2.78e-05
.param mcrdlm2p1_cc_w_1_120_s_3_500=1.13e-11
.param mcrdlm2p1_cf_w_1_120_s_3_500=3.04e-11
.param mcrdlm2l1_ca_w_0_140_s_0_140=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_140=1.03e-10
.param mcrdlm2l1_cf_w_0_140_s_0_140=2.76e-12
.param mcrdlm2l1_ca_w_0_140_s_0_175=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_175=1.01e-10
.param mcrdlm2l1_cf_w_0_140_s_0_175=3.45e-12
.param mcrdlm2l1_ca_w_0_140_s_0_210=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_210=9.59e-11
.param mcrdlm2l1_cf_w_0_140_s_0_210=4.15e-12
.param mcrdlm2l1_ca_w_0_140_s_0_280=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_280=8.47e-11
.param mcrdlm2l1_cf_w_0_140_s_0_280=5.51e-12
.param mcrdlm2l1_ca_w_0_140_s_0_350=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_350=7.32e-11
.param mcrdlm2l1_cf_w_0_140_s_0_350=6.83e-12
.param mcrdlm2l1_ca_w_0_140_s_0_420=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_420=6.35e-11
.param mcrdlm2l1_cf_w_0_140_s_0_420=8.16e-12
.param mcrdlm2l1_ca_w_0_140_s_0_560=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_560=5.06e-11
.param mcrdlm2l1_cf_w_0_140_s_0_560=1.06e-11
.param mcrdlm2l1_ca_w_0_140_s_0_840=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_0_840=3.58e-11
.param mcrdlm2l1_cf_w_0_140_s_0_840=1.51e-11
.param mcrdlm2l1_ca_w_0_140_s_1_540=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_1_540=1.95e-11
.param mcrdlm2l1_cf_w_0_140_s_1_540=2.37e-11
.param mcrdlm2l1_ca_w_0_140_s_3_500=4.01e-05
.param mcrdlm2l1_cc_w_0_140_s_3_500=5.89e-12
.param mcrdlm2l1_cf_w_0_140_s_3_500=3.47e-11
.param mcrdlm2l1_ca_w_1_120_s_0_140=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_140=1.24e-10
.param mcrdlm2l1_cf_w_1_120_s_0_140=2.80e-12
.param mcrdlm2l1_ca_w_1_120_s_0_175=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_175=1.21e-10
.param mcrdlm2l1_cf_w_1_120_s_0_175=3.50e-12
.param mcrdlm2l1_ca_w_1_120_s_0_210=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_210=1.15e-10
.param mcrdlm2l1_cf_w_1_120_s_0_210=4.19e-12
.param mcrdlm2l1_ca_w_1_120_s_0_280=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_280=1.01e-10
.param mcrdlm2l1_cf_w_1_120_s_0_280=5.55e-12
.param mcrdlm2l1_ca_w_1_120_s_0_350=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_350=8.78e-11
.param mcrdlm2l1_cf_w_1_120_s_0_350=6.88e-12
.param mcrdlm2l1_ca_w_1_120_s_0_420=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_420=7.71e-11
.param mcrdlm2l1_cf_w_1_120_s_0_420=8.17e-12
.param mcrdlm2l1_ca_w_1_120_s_0_560=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_560=6.20e-11
.param mcrdlm2l1_cf_w_1_120_s_0_560=1.07e-11
.param mcrdlm2l1_ca_w_1_120_s_0_840=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_0_840=4.49e-11
.param mcrdlm2l1_cf_w_1_120_s_0_840=1.52e-11
.param mcrdlm2l1_ca_w_1_120_s_1_540=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_1_540=2.57e-11
.param mcrdlm2l1_cf_w_1_120_s_1_540=2.43e-11
.param mcrdlm2l1_ca_w_1_120_s_3_500=4.01e-05
.param mcrdlm2l1_cc_w_1_120_s_3_500=8.76e-12
.param mcrdlm2l1_cf_w_1_120_s_3_500=3.70e-11
.param mcrdlm2m1_ca_w_0_140_s_0_140=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_140=9.48e-11
.param mcrdlm2m1_cf_w_0_140_s_0_140=8.45e-12
.param mcrdlm2m1_ca_w_0_140_s_0_175=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_175=9.20e-11
.param mcrdlm2m1_cf_w_0_140_s_0_175=1.07e-11
.param mcrdlm2m1_ca_w_0_140_s_0_210=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_210=8.60e-11
.param mcrdlm2m1_cf_w_0_140_s_0_210=1.29e-11
.param mcrdlm2m1_ca_w_0_140_s_0_280=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_280=7.41e-11
.param mcrdlm2m1_cf_w_0_140_s_0_280=1.69e-11
.param mcrdlm2m1_ca_w_0_140_s_0_350=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_350=6.26e-11
.param mcrdlm2m1_cf_w_0_140_s_0_350=2.06e-11
.param mcrdlm2m1_ca_w_0_140_s_0_420=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_420=5.25e-11
.param mcrdlm2m1_cf_w_0_140_s_0_420=2.40e-11
.param mcrdlm2m1_ca_w_0_140_s_0_560=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_560=3.93e-11
.param mcrdlm2m1_cf_w_0_140_s_0_560=3.00e-11
.param mcrdlm2m1_ca_w_0_140_s_0_840=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_0_840=2.49e-11
.param mcrdlm2m1_cf_w_0_140_s_0_840=3.87e-11
.param mcrdlm2m1_ca_w_0_140_s_1_540=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_1_540=1.08e-11
.param mcrdlm2m1_cf_w_0_140_s_1_540=5.05e-11
.param mcrdlm2m1_ca_w_0_140_s_3_500=1.31e-04
.param mcrdlm2m1_cc_w_0_140_s_3_500=2.50e-12
.param mcrdlm2m1_cf_w_0_140_s_3_500=5.87e-11
.param mcrdlm2m1_ca_w_1_120_s_0_140=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_140=1.11e-10
.param mcrdlm2m1_cf_w_1_120_s_0_140=8.46e-12
.param mcrdlm2m1_ca_w_1_120_s_0_175=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_175=1.08e-10
.param mcrdlm2m1_cf_w_1_120_s_0_175=1.07e-11
.param mcrdlm2m1_ca_w_1_120_s_0_210=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_210=1.02e-10
.param mcrdlm2m1_cf_w_1_120_s_0_210=1.29e-11
.param mcrdlm2m1_ca_w_1_120_s_0_280=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_280=8.75e-11
.param mcrdlm2m1_cf_w_1_120_s_0_280=1.69e-11
.param mcrdlm2m1_ca_w_1_120_s_0_350=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_350=7.44e-11
.param mcrdlm2m1_cf_w_1_120_s_0_350=2.07e-11
.param mcrdlm2m1_ca_w_1_120_s_0_420=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_420=6.42e-11
.param mcrdlm2m1_cf_w_1_120_s_0_420=2.40e-11
.param mcrdlm2m1_ca_w_1_120_s_0_560=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_560=4.93e-11
.param mcrdlm2m1_cf_w_1_120_s_0_560=2.99e-11
.param mcrdlm2m1_ca_w_1_120_s_0_840=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_0_840=3.31e-11
.param mcrdlm2m1_cf_w_1_120_s_0_840=3.90e-11
.param mcrdlm2m1_ca_w_1_120_s_1_540=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_1_540=1.65e-11
.param mcrdlm2m1_cf_w_1_120_s_1_540=5.16e-11
.param mcrdlm2m1_ca_w_1_120_s_3_500=1.31e-04
.param mcrdlm2m1_cc_w_1_120_s_3_500=4.73e-12
.param mcrdlm2m1_cf_w_1_120_s_3_500=6.29e-11
.param mcm4m3f_ca_w_0_300_s_0_300=1.01e-04
.param mcm4m3f_cc_w_0_300_s_0_300=9.07e-11
.param mcm4m3f_cf_w_0_300_s_0_300=1.28e-11
.param mcm4m3f_ca_w_0_300_s_0_360=1.01e-04
.param mcm4m3f_cc_w_0_300_s_0_360=8.30e-11
.param mcm4m3f_cf_w_0_300_s_0_360=1.51e-11
.param mcm4m3f_ca_w_0_300_s_0_450=1.01e-04
.param mcm4m3f_cc_w_0_300_s_0_450=7.20e-11
.param mcm4m3f_cf_w_0_300_s_0_450=1.84e-11
.param mcm4m3f_ca_w_0_300_s_0_600=1.01e-04
.param mcm4m3f_cc_w_0_300_s_0_600=5.84e-11
.param mcm4m3f_cf_w_0_300_s_0_600=2.34e-11
.param mcm4m3f_ca_w_0_300_s_0_800=1.01e-04
.param mcm4m3f_cc_w_0_300_s_0_800=4.47e-11
.param mcm4m3f_cf_w_0_300_s_0_800=2.91e-11
.param mcm4m3f_ca_w_0_300_s_1_000=1.01e-04
.param mcm4m3f_cc_w_0_300_s_1_000=3.47e-11
.param mcm4m3f_cf_w_0_300_s_1_000=3.40e-11
.param mcm4m3f_ca_w_0_300_s_1_200=1.01e-04
.param mcm4m3f_cc_w_0_300_s_1_200=2.74e-11
.param mcm4m3f_cf_w_0_300_s_1_200=3.81e-11
.param mcm4m3f_ca_w_0_300_s_2_100=1.01e-04
.param mcm4m3f_cc_w_0_300_s_2_100=1.09e-11
.param mcm4m3f_cf_w_0_300_s_2_100=4.98e-11
.param mcm4m3f_ca_w_0_300_s_3_300=1.01e-04
.param mcm4m3f_cc_w_0_300_s_3_300=3.74e-12
.param mcm4m3f_cf_w_0_300_s_3_300=5.62e-11
.param mcm4m3f_ca_w_0_300_s_9_000=1.01e-04
.param mcm4m3f_cc_w_0_300_s_9_000=1.10e-13
.param mcm4m3f_cf_w_0_300_s_9_000=5.97e-11
.param mcm4m3f_ca_w_2_400_s_0_300=1.01e-04
.param mcm4m3f_cc_w_2_400_s_0_300=9.86e-11
.param mcm4m3f_cf_w_2_400_s_0_300=1.29e-11
.param mcm4m3f_ca_w_2_400_s_0_360=1.01e-04
.param mcm4m3f_cc_w_2_400_s_0_360=9.03e-11
.param mcm4m3f_cf_w_2_400_s_0_360=1.52e-11
.param mcm4m3f_ca_w_2_400_s_0_450=1.01e-04
.param mcm4m3f_cc_w_2_400_s_0_450=7.89e-11
.param mcm4m3f_cf_w_2_400_s_0_450=1.84e-11
.param mcm4m3f_ca_w_2_400_s_0_600=1.01e-04
.param mcm4m3f_cc_w_2_400_s_0_600=6.39e-11
.param mcm4m3f_cf_w_2_400_s_0_600=2.34e-11
.param mcm4m3f_ca_w_2_400_s_0_800=1.01e-04
.param mcm4m3f_cc_w_2_400_s_0_800=4.92e-11
.param mcm4m3f_cf_w_2_400_s_0_800=2.92e-11
.param mcm4m3f_ca_w_2_400_s_1_000=1.01e-04
.param mcm4m3f_cc_w_2_400_s_1_000=3.85e-11
.param mcm4m3f_cf_w_2_400_s_1_000=3.42e-11
.param mcm4m3f_ca_w_2_400_s_1_200=1.01e-04
.param mcm4m3f_cc_w_2_400_s_1_200=3.07e-11
.param mcm4m3f_cf_w_2_400_s_1_200=3.83e-11
.param mcm4m3f_ca_w_2_400_s_2_100=1.01e-04
.param mcm4m3f_cc_w_2_400_s_2_100=1.27e-11
.param mcm4m3f_cf_w_2_400_s_2_100=5.06e-11
.param mcm4m3f_ca_w_2_400_s_3_300=1.01e-04
.param mcm4m3f_cc_w_2_400_s_3_300=4.61e-12
.param mcm4m3f_cf_w_2_400_s_3_300=5.78e-11
.param mcm4m3f_ca_w_2_400_s_9_000=1.01e-04
.param mcm4m3f_cc_w_2_400_s_9_000=1.40e-13
.param mcm4m3f_cf_w_2_400_s_9_000=6.21e-11
.param mcm4m3d_ca_w_0_300_s_0_300=1.03e-04
.param mcm4m3d_cc_w_0_300_s_0_300=9.03e-11
.param mcm4m3d_cf_w_0_300_s_0_300=1.30e-11
.param mcm4m3d_ca_w_0_300_s_0_360=1.03e-04
.param mcm4m3d_cc_w_0_300_s_0_360=8.26e-11
.param mcm4m3d_cf_w_0_300_s_0_360=1.54e-11
.param mcm4m3d_ca_w_0_300_s_0_450=1.03e-04
.param mcm4m3d_cc_w_0_300_s_0_450=7.16e-11
.param mcm4m3d_cf_w_0_300_s_0_450=1.87e-11
.param mcm4m3d_ca_w_0_300_s_0_600=1.03e-04
.param mcm4m3d_cc_w_0_300_s_0_600=5.79e-11
.param mcm4m3d_cf_w_0_300_s_0_600=2.38e-11
.param mcm4m3d_ca_w_0_300_s_0_800=1.03e-04
.param mcm4m3d_cc_w_0_300_s_0_800=4.41e-11
.param mcm4m3d_cf_w_0_300_s_0_800=2.96e-11
.param mcm4m3d_ca_w_0_300_s_1_000=1.03e-04
.param mcm4m3d_cc_w_0_300_s_1_000=3.41e-11
.param mcm4m3d_cf_w_0_300_s_1_000=3.47e-11
.param mcm4m3d_ca_w_0_300_s_1_200=1.03e-04
.param mcm4m3d_cc_w_0_300_s_1_200=2.68e-11
.param mcm4m3d_cf_w_0_300_s_1_200=3.88e-11
.param mcm4m3d_ca_w_0_300_s_2_100=1.03e-04
.param mcm4m3d_cc_w_0_300_s_2_100=1.03e-11
.param mcm4m3d_cf_w_0_300_s_2_100=5.07e-11
.param mcm4m3d_ca_w_0_300_s_3_300=1.03e-04
.param mcm4m3d_cc_w_0_300_s_3_300=3.34e-12
.param mcm4m3d_cf_w_0_300_s_3_300=5.69e-11
.param mcm4m3d_ca_w_0_300_s_9_000=1.03e-04
.param mcm4m3d_cc_w_0_300_s_9_000=3.00e-14
.param mcm4m3d_cf_w_0_300_s_9_000=6.01e-11
.param mcm4m3d_ca_w_2_400_s_0_300=1.03e-04
.param mcm4m3d_cc_w_2_400_s_0_300=9.75e-11
.param mcm4m3d_cf_w_2_400_s_0_300=1.31e-11
.param mcm4m3d_ca_w_2_400_s_0_360=1.03e-04
.param mcm4m3d_cc_w_2_400_s_0_360=8.91e-11
.param mcm4m3d_cf_w_2_400_s_0_360=1.54e-11
.param mcm4m3d_ca_w_2_400_s_0_450=1.03e-04
.param mcm4m3d_cc_w_2_400_s_0_450=7.76e-11
.param mcm4m3d_cf_w_2_400_s_0_450=1.88e-11
.param mcm4m3d_ca_w_2_400_s_0_600=1.03e-04
.param mcm4m3d_cc_w_2_400_s_0_600=6.27e-11
.param mcm4m3d_cf_w_2_400_s_0_600=2.39e-11
.param mcm4m3d_ca_w_2_400_s_0_800=1.03e-04
.param mcm4m3d_cc_w_2_400_s_0_800=4.80e-11
.param mcm4m3d_cf_w_2_400_s_0_800=2.98e-11
.param mcm4m3d_ca_w_2_400_s_1_000=1.03e-04
.param mcm4m3d_cc_w_2_400_s_1_000=3.73e-11
.param mcm4m3d_cf_w_2_400_s_1_000=3.49e-11
.param mcm4m3d_ca_w_2_400_s_1_200=1.03e-04
.param mcm4m3d_cc_w_2_400_s_1_200=2.95e-11
.param mcm4m3d_cf_w_2_400_s_1_200=3.91e-11
.param mcm4m3d_ca_w_2_400_s_2_100=1.03e-04
.param mcm4m3d_cc_w_2_400_s_2_100=1.18e-11
.param mcm4m3d_cf_w_2_400_s_2_100=5.14e-11
.param mcm4m3d_ca_w_2_400_s_3_300=1.03e-04
.param mcm4m3d_cc_w_2_400_s_3_300=4.00e-12
.param mcm4m3d_cf_w_2_400_s_3_300=5.84e-11
.param mcm4m3d_ca_w_2_400_s_9_000=1.03e-04
.param mcm4m3d_cc_w_2_400_s_9_000=3.50e-14
.param mcm4m3d_cf_w_2_400_s_9_000=6.22e-11
.param mcm4m3p1_ca_w_0_300_s_0_300=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_0_300=8.99e-11
.param mcm4m3p1_cf_w_0_300_s_0_300=1.33e-11
.param mcm4m3p1_ca_w_0_300_s_0_360=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_0_360=8.20e-11
.param mcm4m3p1_cf_w_0_300_s_0_360=1.56e-11
.param mcm4m3p1_ca_w_0_300_s_0_450=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_0_450=7.10e-11
.param mcm4m3p1_cf_w_0_300_s_0_450=1.91e-11
.param mcm4m3p1_ca_w_0_300_s_0_600=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_0_600=5.73e-11
.param mcm4m3p1_cf_w_0_300_s_0_600=2.43e-11
.param mcm4m3p1_ca_w_0_300_s_0_800=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_0_800=4.35e-11
.param mcm4m3p1_cf_w_0_300_s_0_800=3.02e-11
.param mcm4m3p1_ca_w_0_300_s_1_000=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_1_000=3.33e-11
.param mcm4m3p1_cf_w_0_300_s_1_000=3.53e-11
.param mcm4m3p1_ca_w_0_300_s_1_200=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_1_200=2.60e-11
.param mcm4m3p1_cf_w_0_300_s_1_200=3.96e-11
.param mcm4m3p1_ca_w_0_300_s_2_100=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_2_100=9.64e-12
.param mcm4m3p1_cf_w_0_300_s_2_100=5.15e-11
.param mcm4m3p1_ca_w_0_300_s_3_300=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_3_300=2.96e-12
.param mcm4m3p1_cf_w_0_300_s_3_300=5.75e-11
.param mcm4m3p1_ca_w_0_300_s_9_000=1.04e-04
.param mcm4m3p1_cc_w_0_300_s_9_000=3.50e-14
.param mcm4m3p1_cf_w_0_300_s_9_000=6.04e-11
.param mcm4m3p1_ca_w_2_400_s_0_300=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_0_300=9.64e-11
.param mcm4m3p1_cf_w_2_400_s_0_300=1.34e-11
.param mcm4m3p1_ca_w_2_400_s_0_360=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_0_360=8.78e-11
.param mcm4m3p1_cf_w_2_400_s_0_360=1.58e-11
.param mcm4m3p1_ca_w_2_400_s_0_450=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_0_450=7.65e-11
.param mcm4m3p1_cf_w_2_400_s_0_450=1.92e-11
.param mcm4m3p1_ca_w_2_400_s_0_600=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_0_600=6.16e-11
.param mcm4m3p1_cf_w_2_400_s_0_600=2.44e-11
.param mcm4m3p1_ca_w_2_400_s_0_800=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_0_800=4.69e-11
.param mcm4m3p1_cf_w_2_400_s_0_800=3.04e-11
.param mcm4m3p1_ca_w_2_400_s_1_000=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_1_000=3.62e-11
.param mcm4m3p1_cf_w_2_400_s_1_000=3.56e-11
.param mcm4m3p1_ca_w_2_400_s_1_200=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_1_200=2.83e-11
.param mcm4m3p1_cf_w_2_400_s_1_200=3.99e-11
.param mcm4m3p1_ca_w_2_400_s_2_100=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_2_100=1.09e-11
.param mcm4m3p1_cf_w_2_400_s_2_100=5.23e-11
.param mcm4m3p1_ca_w_2_400_s_3_300=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_3_300=3.43e-12
.param mcm4m3p1_cf_w_2_400_s_3_300=5.89e-11
.param mcm4m3p1_ca_w_2_400_s_9_000=1.04e-04
.param mcm4m3p1_cc_w_2_400_s_9_000=4.00e-14
.param mcm4m3p1_cf_w_2_400_s_9_000=6.23e-11
.param mcm4m3l1_ca_w_0_300_s_0_300=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_0_300=8.88e-11
.param mcm4m3l1_cf_w_0_300_s_0_300=1.39e-11
.param mcm4m3l1_ca_w_0_300_s_0_360=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_0_360=8.08e-11
.param mcm4m3l1_cf_w_0_300_s_0_360=1.64e-11
.param mcm4m3l1_ca_w_0_300_s_0_450=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_0_450=7.02e-11
.param mcm4m3l1_cf_w_0_300_s_0_450=2.00e-11
.param mcm4m3l1_ca_w_0_300_s_0_600=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_0_600=5.59e-11
.param mcm4m3l1_cf_w_0_300_s_0_600=2.54e-11
.param mcm4m3l1_ca_w_0_300_s_0_800=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_0_800=4.19e-11
.param mcm4m3l1_cf_w_0_300_s_0_800=3.17e-11
.param mcm4m3l1_ca_w_0_300_s_1_000=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_1_000=3.17e-11
.param mcm4m3l1_cf_w_0_300_s_1_000=3.70e-11
.param mcm4m3l1_ca_w_0_300_s_1_200=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_1_200=2.43e-11
.param mcm4m3l1_cf_w_0_300_s_1_200=4.14e-11
.param mcm4m3l1_ca_w_0_300_s_2_100=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_2_100=8.33e-12
.param mcm4m3l1_cf_w_0_300_s_2_100=5.35e-11
.param mcm4m3l1_ca_w_0_300_s_3_300=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_3_300=2.24e-12
.param mcm4m3l1_cf_w_0_300_s_3_300=5.90e-11
.param mcm4m3l1_ca_w_0_300_s_9_000=1.09e-04
.param mcm4m3l1_cc_w_0_300_s_9_000=5.00e-15
.param mcm4m3l1_cf_w_0_300_s_9_000=6.13e-11
.param mcm4m3l1_ca_w_2_400_s_0_300=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_0_300=9.39e-11
.param mcm4m3l1_cf_w_2_400_s_0_300=1.39e-11
.param mcm4m3l1_ca_w_2_400_s_0_360=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_0_360=8.52e-11
.param mcm4m3l1_cf_w_2_400_s_0_360=1.64e-11
.param mcm4m3l1_ca_w_2_400_s_0_450=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_0_450=7.39e-11
.param mcm4m3l1_cf_w_2_400_s_0_450=2.00e-11
.param mcm4m3l1_ca_w_2_400_s_0_600=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_0_600=5.91e-11
.param mcm4m3l1_cf_w_2_400_s_0_600=2.55e-11
.param mcm4m3l1_ca_w_2_400_s_0_800=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_0_800=4.43e-11
.param mcm4m3l1_cf_w_2_400_s_0_800=3.19e-11
.param mcm4m3l1_ca_w_2_400_s_1_000=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_1_000=3.37e-11
.param mcm4m3l1_cf_w_2_400_s_1_000=3.73e-11
.param mcm4m3l1_ca_w_2_400_s_1_200=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_1_200=2.60e-11
.param mcm4m3l1_cf_w_2_400_s_1_200=4.17e-11
.param mcm4m3l1_ca_w_2_400_s_2_100=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_2_100=9.09e-12
.param mcm4m3l1_cf_w_2_400_s_2_100=5.42e-11
.param mcm4m3l1_ca_w_2_400_s_3_300=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_3_300=2.50e-12
.param mcm4m3l1_cf_w_2_400_s_3_300=6.03e-11
.param mcm4m3l1_ca_w_2_400_s_9_000=1.09e-04
.param mcm4m3l1_cc_w_2_400_s_9_000=0.00e+00
.param mcm4m3l1_cf_w_2_400_s_9_000=6.27e-11
.param mcm4m3m1_ca_w_0_300_s_0_300=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_0_300=8.60e-11
.param mcm4m3m1_cf_w_0_300_s_0_300=1.56e-11
.param mcm4m3m1_ca_w_0_300_s_0_360=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_0_360=7.78e-11
.param mcm4m3m1_cf_w_0_300_s_0_360=1.85e-11
.param mcm4m3m1_ca_w_0_300_s_0_450=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_0_450=6.70e-11
.param mcm4m3m1_cf_w_0_300_s_0_450=2.25e-11
.param mcm4m3m1_ca_w_0_300_s_0_600=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_0_600=5.24e-11
.param mcm4m3m1_cf_w_0_300_s_0_600=2.86e-11
.param mcm4m3m1_ca_w_0_300_s_0_800=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_0_800=3.81e-11
.param mcm4m3m1_cf_w_0_300_s_0_800=3.57e-11
.param mcm4m3m1_ca_w_0_300_s_1_000=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_1_000=2.80e-11
.param mcm4m3m1_cf_w_0_300_s_1_000=4.16e-11
.param mcm4m3m1_ca_w_0_300_s_1_200=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_1_200=2.06e-11
.param mcm4m3m1_cf_w_0_300_s_1_200=4.64e-11
.param mcm4m3m1_ca_w_0_300_s_2_100=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_2_100=5.72e-12
.param mcm4m3m1_cf_w_0_300_s_2_100=5.84e-11
.param mcm4m3m1_ca_w_0_300_s_3_300=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_3_300=1.13e-12
.param mcm4m3m1_cf_w_0_300_s_3_300=6.27e-11
.param mcm4m3m1_ca_w_0_300_s_9_000=1.21e-04
.param mcm4m3m1_cc_w_0_300_s_9_000=3.50e-14
.param mcm4m3m1_cf_w_0_300_s_9_000=6.39e-11
.param mcm4m3m1_ca_w_2_400_s_0_300=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_0_300=8.85e-11
.param mcm4m3m1_cf_w_2_400_s_0_300=1.57e-11
.param mcm4m3m1_ca_w_2_400_s_0_360=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_0_360=7.98e-11
.param mcm4m3m1_cf_w_2_400_s_0_360=1.86e-11
.param mcm4m3m1_ca_w_2_400_s_0_450=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_0_450=6.87e-11
.param mcm4m3m1_cf_w_2_400_s_0_450=2.26e-11
.param mcm4m3m1_ca_w_2_400_s_0_600=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_0_600=5.38e-11
.param mcm4m3m1_cf_w_2_400_s_0_600=2.87e-11
.param mcm4m3m1_ca_w_2_400_s_0_800=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_0_800=3.91e-11
.param mcm4m3m1_cf_w_2_400_s_0_800=3.59e-11
.param mcm4m3m1_ca_w_2_400_s_1_000=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_1_000=2.86e-11
.param mcm4m3m1_cf_w_2_400_s_1_000=4.18e-11
.param mcm4m3m1_ca_w_2_400_s_1_200=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_1_200=2.13e-11
.param mcm4m3m1_cf_w_2_400_s_1_200=4.68e-11
.param mcm4m3m1_ca_w_2_400_s_2_100=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_2_100=5.90e-12
.param mcm4m3m1_cf_w_2_400_s_2_100=5.90e-11
.param mcm4m3m1_ca_w_2_400_s_3_300=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_3_300=1.20e-12
.param mcm4m3m1_cf_w_2_400_s_3_300=6.35e-11
.param mcm4m3m1_ca_w_2_400_s_9_000=1.21e-04
.param mcm4m3m1_cc_w_2_400_s_9_000=5.00e-14
.param mcm4m3m1_cf_w_2_400_s_9_000=6.47e-11
.param mcm4m3m2_ca_w_0_300_s_0_300=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_0_300=7.80e-11
.param mcm4m3m2_cf_w_0_300_s_0_300=2.20e-11
.param mcm4m3m2_ca_w_0_300_s_0_360=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_0_360=6.98e-11
.param mcm4m3m2_cf_w_0_300_s_0_360=2.58e-11
.param mcm4m3m2_ca_w_0_300_s_0_450=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_0_450=5.89e-11
.param mcm4m3m2_cf_w_0_300_s_0_450=3.13e-11
.param mcm4m3m2_ca_w_0_300_s_0_600=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_0_600=4.42e-11
.param mcm4m3m2_cf_w_0_300_s_0_600=3.94e-11
.param mcm4m3m2_ca_w_0_300_s_0_800=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_0_800=3.01e-11
.param mcm4m3m2_cf_w_0_300_s_0_800=4.83e-11
.param mcm4m3m2_ca_w_0_300_s_1_000=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_1_000=2.03e-11
.param mcm4m3m2_cf_w_0_300_s_1_000=5.54e-11
.param mcm4m3m2_ca_w_0_300_s_1_200=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_1_200=1.37e-11
.param mcm4m3m2_cf_w_0_300_s_1_200=6.05e-11
.param mcm4m3m2_ca_w_0_300_s_2_100=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_2_100=2.53e-12
.param mcm4m3m2_cf_w_0_300_s_2_100=7.07e-11
.param mcm4m3m2_ca_w_0_300_s_3_300=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_3_300=3.70e-13
.param mcm4m3m2_cf_w_0_300_s_3_300=7.29e-11
.param mcm4m3m2_ca_w_0_300_s_9_000=1.71e-04
.param mcm4m3m2_cc_w_0_300_s_9_000=2.50e-14
.param mcm4m3m2_cf_w_0_300_s_9_000=7.35e-11
.param mcm4m3m2_ca_w_2_400_s_0_300=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_0_300=7.87e-11
.param mcm4m3m2_cf_w_2_400_s_0_300=2.21e-11
.param mcm4m3m2_ca_w_2_400_s_0_360=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_0_360=7.04e-11
.param mcm4m3m2_cf_w_2_400_s_0_360=2.60e-11
.param mcm4m3m2_ca_w_2_400_s_0_450=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_0_450=5.91e-11
.param mcm4m3m2_cf_w_2_400_s_0_450=3.14e-11
.param mcm4m3m2_ca_w_2_400_s_0_600=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_0_600=4.46e-11
.param mcm4m3m2_cf_w_2_400_s_0_600=3.95e-11
.param mcm4m3m2_ca_w_2_400_s_0_800=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_0_800=3.03e-11
.param mcm4m3m2_cf_w_2_400_s_0_800=4.85e-11
.param mcm4m3m2_ca_w_2_400_s_1_000=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_1_000=2.08e-11
.param mcm4m3m2_cf_w_2_400_s_1_000=5.54e-11
.param mcm4m3m2_ca_w_2_400_s_1_200=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_1_200=1.39e-11
.param mcm4m3m2_cf_w_2_400_s_1_200=6.06e-11
.param mcm4m3m2_ca_w_2_400_s_2_100=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_2_100=2.55e-12
.param mcm4m3m2_cf_w_2_400_s_2_100=7.12e-11
.param mcm4m3m2_ca_w_2_400_s_3_300=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_3_300=3.50e-13
.param mcm4m3m2_cf_w_2_400_s_3_300=7.32e-11
.param mcm4m3m2_ca_w_2_400_s_9_000=1.71e-04
.param mcm4m3m2_cc_w_2_400_s_9_000=5.00e-14
.param mcm4m3m2_cf_w_2_400_s_9_000=7.38e-11
.param mcm5m3f_ca_w_0_300_s_0_300=3.24e-05
.param mcm5m3f_cc_w_0_300_s_0_300=1.02e-10
.param mcm5m3f_cf_w_0_300_s_0_300=4.70e-12
.param mcm5m3f_ca_w_0_300_s_0_360=3.24e-05
.param mcm5m3f_cc_w_0_300_s_0_360=9.41e-11
.param mcm5m3f_cf_w_0_300_s_0_360=5.63e-12
.param mcm5m3f_ca_w_0_300_s_0_450=3.24e-05
.param mcm5m3f_cc_w_0_300_s_0_450=8.44e-11
.param mcm5m3f_cf_w_0_300_s_0_450=7.03e-12
.param mcm5m3f_ca_w_0_300_s_0_600=3.24e-05
.param mcm5m3f_cc_w_0_300_s_0_600=7.08e-11
.param mcm5m3f_cf_w_0_300_s_0_600=9.28e-12
.param mcm5m3f_ca_w_0_300_s_0_800=3.24e-05
.param mcm5m3f_cc_w_0_300_s_0_800=5.71e-11
.param mcm5m3f_cf_w_0_300_s_0_800=1.20e-11
.param mcm5m3f_ca_w_0_300_s_1_000=3.24e-05
.param mcm5m3f_cc_w_0_300_s_1_000=4.70e-11
.param mcm5m3f_cf_w_0_300_s_1_000=1.47e-11
.param mcm5m3f_ca_w_0_300_s_1_200=3.24e-05
.param mcm5m3f_cc_w_0_300_s_1_200=3.92e-11
.param mcm5m3f_cf_w_0_300_s_1_200=1.73e-11
.param mcm5m3f_ca_w_0_300_s_2_100=3.24e-05
.param mcm5m3f_cc_w_0_300_s_2_100=2.02e-11
.param mcm5m3f_cf_w_0_300_s_2_100=2.66e-11
.param mcm5m3f_ca_w_0_300_s_3_300=3.24e-05
.param mcm5m3f_cc_w_0_300_s_3_300=9.34e-12
.param mcm5m3f_cf_w_0_300_s_3_300=3.43e-11
.param mcm5m3f_ca_w_0_300_s_9_000=3.24e-05
.param mcm5m3f_cc_w_0_300_s_9_000=3.50e-13
.param mcm5m3f_cf_w_0_300_s_9_000=4.24e-11
.param mcm5m3f_ca_w_2_400_s_0_300=3.24e-05
.param mcm5m3f_cc_w_2_400_s_0_300=1.14e-10
.param mcm5m3f_cf_w_2_400_s_0_300=4.75e-12
.param mcm5m3f_ca_w_2_400_s_0_360=3.24e-05
.param mcm5m3f_cc_w_2_400_s_0_360=1.06e-10
.param mcm5m3f_cf_w_2_400_s_0_360=5.67e-12
.param mcm5m3f_ca_w_2_400_s_0_450=3.24e-05
.param mcm5m3f_cc_w_2_400_s_0_450=9.43e-11
.param mcm5m3f_cf_w_2_400_s_0_450=7.03e-12
.param mcm5m3f_ca_w_2_400_s_0_600=3.24e-05
.param mcm5m3f_cc_w_2_400_s_0_600=7.93e-11
.param mcm5m3f_cf_w_2_400_s_0_600=9.27e-12
.param mcm5m3f_ca_w_2_400_s_0_800=3.24e-05
.param mcm5m3f_cc_w_2_400_s_0_800=6.40e-11
.param mcm5m3f_cf_w_2_400_s_0_800=1.21e-11
.param mcm5m3f_ca_w_2_400_s_1_000=3.24e-05
.param mcm5m3f_cc_w_2_400_s_1_000=5.27e-11
.param mcm5m3f_cf_w_2_400_s_1_000=1.49e-11
.param mcm5m3f_ca_w_2_400_s_1_200=3.24e-05
.param mcm5m3f_cc_w_2_400_s_1_200=4.42e-11
.param mcm5m3f_cf_w_2_400_s_1_200=1.75e-11
.param mcm5m3f_ca_w_2_400_s_2_100=3.24e-05
.param mcm5m3f_cc_w_2_400_s_2_100=2.29e-11
.param mcm5m3f_cf_w_2_400_s_2_100=2.72e-11
.param mcm5m3f_ca_w_2_400_s_3_300=3.24e-05
.param mcm5m3f_cc_w_2_400_s_3_300=1.08e-11
.param mcm5m3f_cf_w_2_400_s_3_300=3.56e-11
.param mcm5m3f_ca_w_2_400_s_9_000=3.24e-05
.param mcm5m3f_cc_w_2_400_s_9_000=4.15e-13
.param mcm5m3f_cf_w_2_400_s_9_000=4.50e-11
.param mcm5m3d_ca_w_0_300_s_0_300=3.40e-05
.param mcm5m3d_cc_w_0_300_s_0_300=1.01e-10
.param mcm5m3d_cf_w_0_300_s_0_300=4.94e-12
.param mcm5m3d_ca_w_0_300_s_0_360=3.40e-05
.param mcm5m3d_cc_w_0_300_s_0_360=9.37e-11
.param mcm5m3d_cf_w_0_300_s_0_360=5.91e-12
.param mcm5m3d_ca_w_0_300_s_0_450=3.40e-05
.param mcm5m3d_cc_w_0_300_s_0_450=8.39e-11
.param mcm5m3d_cf_w_0_300_s_0_450=7.38e-12
.param mcm5m3d_ca_w_0_300_s_0_600=3.40e-05
.param mcm5m3d_cc_w_0_300_s_0_600=7.03e-11
.param mcm5m3d_cf_w_0_300_s_0_600=9.72e-12
.param mcm5m3d_ca_w_0_300_s_0_800=3.40e-05
.param mcm5m3d_cc_w_0_300_s_0_800=5.64e-11
.param mcm5m3d_cf_w_0_300_s_0_800=1.26e-11
.param mcm5m3d_ca_w_0_300_s_1_000=3.40e-05
.param mcm5m3d_cc_w_0_300_s_1_000=4.64e-11
.param mcm5m3d_cf_w_0_300_s_1_000=1.54e-11
.param mcm5m3d_ca_w_0_300_s_1_200=3.40e-05
.param mcm5m3d_cc_w_0_300_s_1_200=3.85e-11
.param mcm5m3d_cf_w_0_300_s_1_200=1.81e-11
.param mcm5m3d_ca_w_0_300_s_2_100=3.40e-05
.param mcm5m3d_cc_w_0_300_s_2_100=1.94e-11
.param mcm5m3d_cf_w_0_300_s_2_100=2.77e-11
.param mcm5m3d_ca_w_0_300_s_3_300=3.40e-05
.param mcm5m3d_cc_w_0_300_s_3_300=8.69e-12
.param mcm5m3d_cf_w_0_300_s_3_300=3.55e-11
.param mcm5m3d_ca_w_0_300_s_9_000=3.40e-05
.param mcm5m3d_cc_w_0_300_s_9_000=2.80e-13
.param mcm5m3d_cf_w_0_300_s_9_000=4.31e-11
.param mcm5m3d_ca_w_2_400_s_0_300=3.40e-05
.param mcm5m3d_cc_w_2_400_s_0_300=1.13e-10
.param mcm5m3d_cf_w_2_400_s_0_300=4.99e-12
.param mcm5m3d_ca_w_2_400_s_0_360=3.40e-05
.param mcm5m3d_cc_w_2_400_s_0_360=1.05e-10
.param mcm5m3d_cf_w_2_400_s_0_360=5.96e-12
.param mcm5m3d_ca_w_2_400_s_0_450=3.40e-05
.param mcm5m3d_cc_w_2_400_s_0_450=9.32e-11
.param mcm5m3d_cf_w_2_400_s_0_450=7.39e-12
.param mcm5m3d_ca_w_2_400_s_0_600=3.40e-05
.param mcm5m3d_cc_w_2_400_s_0_600=7.81e-11
.param mcm5m3d_cf_w_2_400_s_0_600=9.73e-12
.param mcm5m3d_ca_w_2_400_s_0_800=3.40e-05
.param mcm5m3d_cc_w_2_400_s_0_800=6.28e-11
.param mcm5m3d_cf_w_2_400_s_0_800=1.27e-11
.param mcm5m3d_ca_w_2_400_s_1_000=3.40e-05
.param mcm5m3d_cc_w_2_400_s_1_000=5.15e-11
.param mcm5m3d_cf_w_2_400_s_1_000=1.56e-11
.param mcm5m3d_ca_w_2_400_s_1_200=3.40e-05
.param mcm5m3d_cc_w_2_400_s_1_200=4.30e-11
.param mcm5m3d_cf_w_2_400_s_1_200=1.83e-11
.param mcm5m3d_ca_w_2_400_s_2_100=3.40e-05
.param mcm5m3d_cc_w_2_400_s_2_100=2.18e-11
.param mcm5m3d_cf_w_2_400_s_2_100=2.83e-11
.param mcm5m3d_ca_w_2_400_s_3_300=3.40e-05
.param mcm5m3d_cc_w_2_400_s_3_300=9.86e-12
.param mcm5m3d_cf_w_2_400_s_3_300=3.69e-11
.param mcm5m3d_ca_w_2_400_s_9_000=3.40e-05
.param mcm5m3d_cc_w_2_400_s_9_000=3.20e-13
.param mcm5m3d_cf_w_2_400_s_9_000=4.56e-11
.param mcm5m3p1_ca_w_0_300_s_0_300=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_0_300=1.01e-10
.param mcm5m3p1_cf_w_0_300_s_0_300=5.19e-12
.param mcm5m3p1_ca_w_0_300_s_0_360=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_0_360=9.32e-11
.param mcm5m3p1_cf_w_0_300_s_0_360=6.21e-12
.param mcm5m3p1_ca_w_0_300_s_0_450=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_0_450=8.31e-11
.param mcm5m3p1_cf_w_0_300_s_0_450=7.74e-12
.param mcm5m3p1_ca_w_0_300_s_0_600=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_0_600=6.97e-11
.param mcm5m3p1_cf_w_0_300_s_0_600=1.02e-11
.param mcm5m3p1_ca_w_0_300_s_0_800=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_0_800=5.57e-11
.param mcm5m3p1_cf_w_0_300_s_0_800=1.32e-11
.param mcm5m3p1_ca_w_0_300_s_1_000=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_1_000=4.56e-11
.param mcm5m3p1_cf_w_0_300_s_1_000=1.62e-11
.param mcm5m3p1_ca_w_0_300_s_1_200=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_1_200=3.78e-11
.param mcm5m3p1_cf_w_0_300_s_1_200=1.89e-11
.param mcm5m3p1_ca_w_0_300_s_2_100=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_2_100=1.85e-11
.param mcm5m3p1_cf_w_0_300_s_2_100=2.88e-11
.param mcm5m3p1_ca_w_0_300_s_3_300=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_3_300=8.07e-12
.param mcm5m3p1_cf_w_0_300_s_3_300=3.66e-11
.param mcm5m3p1_ca_w_0_300_s_9_000=3.57e-05
.param mcm5m3p1_cc_w_0_300_s_9_000=2.20e-13
.param mcm5m3p1_cf_w_0_300_s_9_000=4.38e-11
.param mcm5m3p1_ca_w_2_400_s_0_300=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_0_300=1.12e-10
.param mcm5m3p1_cf_w_2_400_s_0_300=5.28e-12
.param mcm5m3p1_ca_w_2_400_s_0_360=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_0_360=1.04e-10
.param mcm5m3p1_cf_w_2_400_s_0_360=6.28e-12
.param mcm5m3p1_ca_w_2_400_s_0_450=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_0_450=9.20e-11
.param mcm5m3p1_cf_w_2_400_s_0_450=7.78e-12
.param mcm5m3p1_ca_w_2_400_s_0_600=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_0_600=7.69e-11
.param mcm5m3p1_cf_w_2_400_s_0_600=1.02e-11
.param mcm5m3p1_ca_w_2_400_s_0_800=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_0_800=6.15e-11
.param mcm5m3p1_cf_w_2_400_s_0_800=1.34e-11
.param mcm5m3p1_ca_w_2_400_s_1_000=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_1_000=5.03e-11
.param mcm5m3p1_cf_w_2_400_s_1_000=1.64e-11
.param mcm5m3p1_ca_w_2_400_s_1_200=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_1_200=4.18e-11
.param mcm5m3p1_cf_w_2_400_s_1_200=1.92e-11
.param mcm5m3p1_ca_w_2_400_s_2_100=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_2_100=2.07e-11
.param mcm5m3p1_cf_w_2_400_s_2_100=2.95e-11
.param mcm5m3p1_ca_w_2_400_s_3_300=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_3_300=9.06e-12
.param mcm5m3p1_cf_w_2_400_s_3_300=3.80e-11
.param mcm5m3p1_ca_w_2_400_s_9_000=3.57e-05
.param mcm5m3p1_cc_w_2_400_s_9_000=2.35e-13
.param mcm5m3p1_cf_w_2_400_s_9_000=4.61e-11
.param mcm5m3l1_ca_w_0_300_s_0_300=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_0_300=9.96e-11
.param mcm5m3l1_cf_w_0_300_s_0_300=5.80e-12
.param mcm5m3l1_ca_w_0_300_s_0_360=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_0_360=9.23e-11
.param mcm5m3l1_cf_w_0_300_s_0_360=6.92e-12
.param mcm5m3l1_ca_w_0_300_s_0_450=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_0_450=8.21e-11
.param mcm5m3l1_cf_w_0_300_s_0_450=8.63e-12
.param mcm5m3l1_ca_w_0_300_s_0_600=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_0_600=6.83e-11
.param mcm5m3l1_cf_w_0_300_s_0_600=1.13e-11
.param mcm5m3l1_ca_w_0_300_s_0_800=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_0_800=5.42e-11
.param mcm5m3l1_cf_w_0_300_s_0_800=1.47e-11
.param mcm5m3l1_ca_w_0_300_s_1_000=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_1_000=4.40e-11
.param mcm5m3l1_cf_w_0_300_s_1_000=1.79e-11
.param mcm5m3l1_ca_w_0_300_s_1_200=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_1_200=3.61e-11
.param mcm5m3l1_cf_w_0_300_s_1_200=2.09e-11
.param mcm5m3l1_ca_w_0_300_s_2_100=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_2_100=1.68e-11
.param mcm5m3l1_cf_w_0_300_s_2_100=3.14e-11
.param mcm5m3l1_ca_w_0_300_s_3_300=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_3_300=6.77e-12
.param mcm5m3l1_cf_w_0_300_s_3_300=3.92e-11
.param mcm5m3l1_ca_w_0_300_s_9_000=4.00e-05
.param mcm5m3l1_cc_w_0_300_s_9_000=1.55e-13
.param mcm5m3l1_cf_w_0_300_s_9_000=4.54e-11
.param mcm5m3l1_ca_w_2_400_s_0_300=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_0_300=1.10e-10
.param mcm5m3l1_cf_w_2_400_s_0_300=5.84e-12
.param mcm5m3l1_ca_w_2_400_s_0_360=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_0_360=1.01e-10
.param mcm5m3l1_cf_w_2_400_s_0_360=6.97e-12
.param mcm5m3l1_ca_w_2_400_s_0_450=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_0_450=8.94e-11
.param mcm5m3l1_cf_w_2_400_s_0_450=8.65e-12
.param mcm5m3l1_ca_w_2_400_s_0_600=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_0_600=7.43e-11
.param mcm5m3l1_cf_w_2_400_s_0_600=1.13e-11
.param mcm5m3l1_ca_w_2_400_s_0_800=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_0_800=5.91e-11
.param mcm5m3l1_cf_w_2_400_s_0_800=1.48e-11
.param mcm5m3l1_ca_w_2_400_s_1_000=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_1_000=4.79e-11
.param mcm5m3l1_cf_w_2_400_s_1_000=1.82e-11
.param mcm5m3l1_ca_w_2_400_s_1_200=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_1_200=3.93e-11
.param mcm5m3l1_cf_w_2_400_s_1_200=2.12e-11
.param mcm5m3l1_ca_w_2_400_s_2_100=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_2_100=1.86e-11
.param mcm5m3l1_cf_w_2_400_s_2_100=3.21e-11
.param mcm5m3l1_ca_w_2_400_s_3_300=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_3_300=7.52e-12
.param mcm5m3l1_cf_w_2_400_s_3_300=4.06e-11
.param mcm5m3l1_ca_w_2_400_s_9_000=4.00e-05
.param mcm5m3l1_cc_w_2_400_s_9_000=1.65e-13
.param mcm5m3l1_cf_w_2_400_s_9_000=4.74e-11
.param mcm5m3m1_ca_w_0_300_s_0_300=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_0_300=9.70e-11
.param mcm5m3m1_cf_w_0_300_s_0_300=7.58e-12
.param mcm5m3m1_ca_w_0_300_s_0_360=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_0_360=8.92e-11
.param mcm5m3m1_cf_w_0_300_s_0_360=9.02e-12
.param mcm5m3m1_ca_w_0_300_s_0_450=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_0_450=7.89e-11
.param mcm5m3m1_cf_w_0_300_s_0_450=1.12e-11
.param mcm5m3m1_ca_w_0_300_s_0_600=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_0_600=6.46e-11
.param mcm5m3m1_cf_w_0_300_s_0_600=1.46e-11
.param mcm5m3m1_ca_w_0_300_s_0_800=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_0_800=5.04e-11
.param mcm5m3m1_cf_w_0_300_s_0_800=1.88e-11
.param mcm5m3m1_ca_w_0_300_s_1_000=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_1_000=3.99e-11
.param mcm5m3m1_cf_w_0_300_s_1_000=2.28e-11
.param mcm5m3m1_ca_w_0_300_s_1_200=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_1_200=3.21e-11
.param mcm5m3m1_cf_w_0_300_s_1_200=2.63e-11
.param mcm5m3m1_ca_w_0_300_s_2_100=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_2_100=1.34e-11
.param mcm5m3m1_cf_w_0_300_s_2_100=3.79e-11
.param mcm5m3m1_ca_w_0_300_s_3_300=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_3_300=4.63e-12
.param mcm5m3m1_cf_w_0_300_s_3_300=4.53e-11
.param mcm5m3m1_ca_w_0_300_s_9_000=5.27e-05
.param mcm5m3m1_cc_w_0_300_s_9_000=7.00e-14
.param mcm5m3m1_cf_w_0_300_s_9_000=4.97e-11
.param mcm5m3m1_ca_w_2_400_s_0_300=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_0_300=1.05e-10
.param mcm5m3m1_cf_w_2_400_s_0_300=7.59e-12
.param mcm5m3m1_ca_w_2_400_s_0_360=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_0_360=9.57e-11
.param mcm5m3m1_cf_w_2_400_s_0_360=9.05e-12
.param mcm5m3m1_ca_w_2_400_s_0_450=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_0_450=8.42e-11
.param mcm5m3m1_cf_w_2_400_s_0_450=1.12e-11
.param mcm5m3m1_ca_w_2_400_s_0_600=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_0_600=6.91e-11
.param mcm5m3m1_cf_w_2_400_s_0_600=1.46e-11
.param mcm5m3m1_ca_w_2_400_s_0_800=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_0_800=5.39e-11
.param mcm5m3m1_cf_w_2_400_s_0_800=1.89e-11
.param mcm5m3m1_ca_w_2_400_s_1_000=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_1_000=4.27e-11
.param mcm5m3m1_cf_w_2_400_s_1_000=2.30e-11
.param mcm5m3m1_ca_w_2_400_s_1_200=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_1_200=3.43e-11
.param mcm5m3m1_cf_w_2_400_s_1_200=2.66e-11
.param mcm5m3m1_ca_w_2_400_s_2_100=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_2_100=1.45e-11
.param mcm5m3m1_cf_w_2_400_s_2_100=3.86e-11
.param mcm5m3m1_ca_w_2_400_s_3_300=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_3_300=5.05e-12
.param mcm5m3m1_cf_w_2_400_s_3_300=4.65e-11
.param mcm5m3m1_ca_w_2_400_s_9_000=5.27e-05
.param mcm5m3m1_cc_w_2_400_s_9_000=8.00e-14
.param mcm5m3m1_cf_w_2_400_s_9_000=5.13e-11
.param mcm5m3m2_ca_w_0_300_s_0_300=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_0_300=8.92e-11
.param mcm5m3m2_cf_w_0_300_s_0_300=1.39e-11
.param mcm5m3m2_ca_w_0_300_s_0_360=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_0_360=8.10e-11
.param mcm5m3m2_cf_w_0_300_s_0_360=1.65e-11
.param mcm5m3m2_ca_w_0_300_s_0_450=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_0_450=7.04e-11
.param mcm5m3m2_cf_w_0_300_s_0_450=2.00e-11
.param mcm5m3m2_ca_w_0_300_s_0_600=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_0_600=5.62e-11
.param mcm5m3m2_cf_w_0_300_s_0_600=2.54e-11
.param mcm5m3m2_ca_w_0_300_s_0_800=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_0_800=4.23e-11
.param mcm5m3m2_cf_w_0_300_s_0_800=3.16e-11
.param mcm5m3m2_ca_w_0_300_s_1_000=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_1_000=3.20e-11
.param mcm5m3m2_cf_w_0_300_s_1_000=3.70e-11
.param mcm5m3m2_ca_w_0_300_s_1_200=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_1_200=2.46e-11
.param mcm5m3m2_cf_w_0_300_s_1_200=4.15e-11
.param mcm5m3m2_ca_w_0_300_s_2_100=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_2_100=8.49e-12
.param mcm5m3m2_cf_w_0_300_s_2_100=5.35e-11
.param mcm5m3m2_ca_w_0_300_s_3_300=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_3_300=2.28e-12
.param mcm5m3m2_cf_w_0_300_s_3_300=5.91e-11
.param mcm5m3m2_ca_w_0_300_s_9_000=1.02e-04
.param mcm5m3m2_cc_w_0_300_s_9_000=5.00e-14
.param mcm5m3m2_cf_w_0_300_s_9_000=6.16e-11
.param mcm5m3m2_ca_w_2_400_s_0_300=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_0_300=9.45e-11
.param mcm5m3m2_cf_w_2_400_s_0_300=1.40e-11
.param mcm5m3m2_ca_w_2_400_s_0_360=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_0_360=8.58e-11
.param mcm5m3m2_cf_w_2_400_s_0_360=1.64e-11
.param mcm5m3m2_ca_w_2_400_s_0_450=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_0_450=7.46e-11
.param mcm5m3m2_cf_w_2_400_s_0_450=2.00e-11
.param mcm5m3m2_ca_w_2_400_s_0_600=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_0_600=5.96e-11
.param mcm5m3m2_cf_w_2_400_s_0_600=2.54e-11
.param mcm5m3m2_ca_w_2_400_s_0_800=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_0_800=4.49e-11
.param mcm5m3m2_cf_w_2_400_s_0_800=3.17e-11
.param mcm5m3m2_ca_w_2_400_s_1_000=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_1_000=3.43e-11
.param mcm5m3m2_cf_w_2_400_s_1_000=3.71e-11
.param mcm5m3m2_ca_w_2_400_s_1_200=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_1_200=2.64e-11
.param mcm5m3m2_cf_w_2_400_s_1_200=4.16e-11
.param mcm5m3m2_ca_w_2_400_s_2_100=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_2_100=9.40e-12
.param mcm5m3m2_cf_w_2_400_s_2_100=5.43e-11
.param mcm5m3m2_ca_w_2_400_s_3_300=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_3_300=2.61e-12
.param mcm5m3m2_cf_w_2_400_s_3_300=6.04e-11
.param mcm5m3m2_ca_w_2_400_s_9_000=1.02e-04
.param mcm5m3m2_cc_w_2_400_s_9_000=1.00e-14
.param mcm5m3m2_cf_w_2_400_s_9_000=6.30e-11
.param mcrdlm3f_ca_w_0_300_s_0_300=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_0_300=1.06e-10
.param mcrdlm3f_cf_w_0_300_s_0_300=2.38e-12
.param mcrdlm3f_ca_w_0_300_s_0_360=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_0_360=9.87e-11
.param mcrdlm3f_cf_w_0_300_s_0_360=2.85e-12
.param mcrdlm3f_ca_w_0_300_s_0_450=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_0_450=8.91e-11
.param mcrdlm3f_cf_w_0_300_s_0_450=3.58e-12
.param mcrdlm3f_ca_w_0_300_s_0_600=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_0_600=7.63e-11
.param mcrdlm3f_cf_w_0_300_s_0_600=4.76e-12
.param mcrdlm3f_ca_w_0_300_s_0_800=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_0_800=6.38e-11
.param mcrdlm3f_cf_w_0_300_s_0_800=6.17e-12
.param mcrdlm3f_ca_w_0_300_s_1_000=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_1_000=5.45e-11
.param mcrdlm3f_cf_w_0_300_s_1_000=7.62e-12
.param mcrdlm3f_ca_w_0_300_s_1_200=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_1_200=4.75e-11
.param mcrdlm3f_cf_w_0_300_s_1_200=9.03e-12
.param mcrdlm3f_ca_w_0_300_s_2_100=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_2_100=2.96e-11
.param mcrdlm3f_cf_w_0_300_s_2_100=1.49e-11
.param mcrdlm3f_ca_w_0_300_s_3_300=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_3_300=1.87e-11
.param mcrdlm3f_cf_w_0_300_s_3_300=2.06e-11
.param mcrdlm3f_ca_w_0_300_s_9_000=1.61e-05
.param mcrdlm3f_cc_w_0_300_s_9_000=3.26e-12
.param mcrdlm3f_cf_w_0_300_s_9_000=3.25e-11
.param mcrdlm3f_ca_w_2_400_s_0_300=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_0_300=1.28e-10
.param mcrdlm3f_cf_w_2_400_s_0_300=2.43e-12
.param mcrdlm3f_ca_w_2_400_s_0_360=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_0_360=1.19e-10
.param mcrdlm3f_cf_w_2_400_s_0_360=2.89e-12
.param mcrdlm3f_ca_w_2_400_s_0_450=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_0_450=1.08e-10
.param mcrdlm3f_cf_w_2_400_s_0_450=3.59e-12
.param mcrdlm3f_ca_w_2_400_s_0_600=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_0_600=9.31e-11
.param mcrdlm3f_cf_w_2_400_s_0_600=4.74e-12
.param mcrdlm3f_ca_w_2_400_s_0_800=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_0_800=7.81e-11
.param mcrdlm3f_cf_w_2_400_s_0_800=6.24e-12
.param mcrdlm3f_ca_w_2_400_s_1_000=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_1_000=6.72e-11
.param mcrdlm3f_cf_w_2_400_s_1_000=7.71e-12
.param mcrdlm3f_ca_w_2_400_s_1_200=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_1_200=5.87e-11
.param mcrdlm3f_cf_w_2_400_s_1_200=9.13e-12
.param mcrdlm3f_ca_w_2_400_s_2_100=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_2_100=3.74e-11
.param mcrdlm3f_cf_w_2_400_s_2_100=1.50e-11
.param mcrdlm3f_ca_w_2_400_s_3_300=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_3_300=2.39e-11
.param mcrdlm3f_cf_w_2_400_s_3_300=2.13e-11
.param mcrdlm3f_ca_w_2_400_s_9_000=1.61e-05
.param mcrdlm3f_cc_w_2_400_s_9_000=4.48e-12
.param mcrdlm3f_cf_w_2_400_s_9_000=3.56e-11
.param mcrdlm3d_ca_w_0_300_s_0_300=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_0_300=1.05e-10
.param mcrdlm3d_cf_w_0_300_s_0_300=2.61e-12
.param mcrdlm3d_ca_w_0_300_s_0_360=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_0_360=9.83e-11
.param mcrdlm3d_cf_w_0_300_s_0_360=3.13e-12
.param mcrdlm3d_ca_w_0_300_s_0_450=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_0_450=8.86e-11
.param mcrdlm3d_cf_w_0_300_s_0_450=3.92e-12
.param mcrdlm3d_ca_w_0_300_s_0_600=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_0_600=7.58e-11
.param mcrdlm3d_cf_w_0_300_s_0_600=5.21e-12
.param mcrdlm3d_ca_w_0_300_s_0_800=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_0_800=6.31e-11
.param mcrdlm3d_cf_w_0_300_s_0_800=6.76e-12
.param mcrdlm3d_ca_w_0_300_s_1_000=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_1_000=5.37e-11
.param mcrdlm3d_cf_w_0_300_s_1_000=8.33e-12
.param mcrdlm3d_ca_w_0_300_s_1_200=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_1_200=4.67e-11
.param mcrdlm3d_cf_w_0_300_s_1_200=9.85e-12
.param mcrdlm3d_ca_w_0_300_s_2_100=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_2_100=2.87e-11
.param mcrdlm3d_cf_w_0_300_s_2_100=1.62e-11
.param mcrdlm3d_ca_w_0_300_s_3_300=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_3_300=1.78e-11
.param mcrdlm3d_cf_w_0_300_s_3_300=2.21e-11
.param mcrdlm3d_ca_w_0_300_s_9_000=1.77e-05
.param mcrdlm3d_cc_w_0_300_s_9_000=2.89e-12
.param mcrdlm3d_cf_w_0_300_s_9_000=3.39e-11
.param mcrdlm3d_ca_w_2_400_s_0_300=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_0_300=1.26e-10
.param mcrdlm3d_cf_w_2_400_s_0_300=2.67e-12
.param mcrdlm3d_ca_w_2_400_s_0_360=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_0_360=1.18e-10
.param mcrdlm3d_cf_w_2_400_s_0_360=3.18e-12
.param mcrdlm3d_ca_w_2_400_s_0_450=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_0_450=1.07e-10
.param mcrdlm3d_cf_w_2_400_s_0_450=3.94e-12
.param mcrdlm3d_ca_w_2_400_s_0_600=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_0_600=9.19e-11
.param mcrdlm3d_cf_w_2_400_s_0_600=5.20e-12
.param mcrdlm3d_ca_w_2_400_s_0_800=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_0_800=7.69e-11
.param mcrdlm3d_cf_w_2_400_s_0_800=6.83e-12
.param mcrdlm3d_ca_w_2_400_s_1_000=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_1_000=6.59e-11
.param mcrdlm3d_cf_w_2_400_s_1_000=8.43e-12
.param mcrdlm3d_ca_w_2_400_s_1_200=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_1_200=5.75e-11
.param mcrdlm3d_cf_w_2_400_s_1_200=9.97e-12
.param mcrdlm3d_ca_w_2_400_s_2_100=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_2_100=3.62e-11
.param mcrdlm3d_cf_w_2_400_s_2_100=1.62e-11
.param mcrdlm3d_ca_w_2_400_s_3_300=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_3_300=2.27e-11
.param mcrdlm3d_cf_w_2_400_s_3_300=2.29e-11
.param mcrdlm3d_ca_w_2_400_s_9_000=1.77e-05
.param mcrdlm3d_cc_w_2_400_s_9_000=4.01e-12
.param mcrdlm3d_cf_w_2_400_s_9_000=3.71e-11
.param mcrdlm3p1_ca_w_0_300_s_0_300=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_0_300=1.05e-10
.param mcrdlm3p1_cf_w_0_300_s_0_300=2.87e-12
.param mcrdlm3p1_ca_w_0_300_s_0_360=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_0_360=9.79e-11
.param mcrdlm3p1_cf_w_0_300_s_0_360=3.43e-12
.param mcrdlm3p1_ca_w_0_300_s_0_450=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_0_450=8.81e-11
.param mcrdlm3p1_cf_w_0_300_s_0_450=4.29e-12
.param mcrdlm3p1_ca_w_0_300_s_0_600=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_0_600=7.51e-11
.param mcrdlm3p1_cf_w_0_300_s_0_600=5.70e-12
.param mcrdlm3p1_ca_w_0_300_s_0_800=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_0_800=6.24e-11
.param mcrdlm3p1_cf_w_0_300_s_0_800=7.37e-12
.param mcrdlm3p1_ca_w_0_300_s_1_000=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_1_000=5.30e-11
.param mcrdlm3p1_cf_w_0_300_s_1_000=9.07e-12
.param mcrdlm3p1_ca_w_0_300_s_1_200=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_1_200=4.59e-11
.param mcrdlm3p1_cf_w_0_300_s_1_200=1.07e-11
.param mcrdlm3p1_ca_w_0_300_s_2_100=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_2_100=2.77e-11
.param mcrdlm3p1_cf_w_0_300_s_2_100=1.74e-11
.param mcrdlm3p1_ca_w_0_300_s_3_300=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_3_300=1.69e-11
.param mcrdlm3p1_cf_w_0_300_s_3_300=2.36e-11
.param mcrdlm3p1_ca_w_0_300_s_9_000=1.94e-05
.param mcrdlm3p1_cc_w_0_300_s_9_000=2.58e-12
.param mcrdlm3p1_cf_w_0_300_s_9_000=3.52e-11
.param mcrdlm3p1_ca_w_2_400_s_0_300=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_0_300=1.25e-10
.param mcrdlm3p1_cf_w_2_400_s_0_300=2.95e-12
.param mcrdlm3p1_ca_w_2_400_s_0_360=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_0_360=1.17e-10
.param mcrdlm3p1_cf_w_2_400_s_0_360=3.50e-12
.param mcrdlm3p1_ca_w_2_400_s_0_450=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_0_450=1.06e-10
.param mcrdlm3p1_cf_w_2_400_s_0_450=4.35e-12
.param mcrdlm3p1_ca_w_2_400_s_0_600=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_0_600=9.07e-11
.param mcrdlm3p1_cf_w_2_400_s_0_600=5.70e-12
.param mcrdlm3p1_ca_w_2_400_s_0_800=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_0_800=7.57e-11
.param mcrdlm3p1_cf_w_2_400_s_0_800=7.48e-12
.param mcrdlm3p1_ca_w_2_400_s_1_000=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_1_000=6.46e-11
.param mcrdlm3p1_cf_w_2_400_s_1_000=9.21e-12
.param mcrdlm3p1_ca_w_2_400_s_1_200=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_1_200=5.62e-11
.param mcrdlm3p1_cf_w_2_400_s_1_200=1.09e-11
.param mcrdlm3p1_ca_w_2_400_s_2_100=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_2_100=3.51e-11
.param mcrdlm3p1_cf_w_2_400_s_2_100=1.75e-11
.param mcrdlm3p1_ca_w_2_400_s_3_300=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_3_300=2.18e-11
.param mcrdlm3p1_cf_w_2_400_s_3_300=2.45e-11
.param mcrdlm3p1_ca_w_2_400_s_9_000=1.94e-05
.param mcrdlm3p1_cc_w_2_400_s_9_000=3.67e-12
.param mcrdlm3p1_cf_w_2_400_s_9_000=3.86e-11
.param mcrdlm3l1_ca_w_0_300_s_0_300=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_0_300=1.04e-10
.param mcrdlm3l1_cf_w_0_300_s_0_300=3.47e-12
.param mcrdlm3l1_ca_w_0_300_s_0_360=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_0_360=9.68e-11
.param mcrdlm3l1_cf_w_0_300_s_0_360=4.15e-12
.param mcrdlm3l1_ca_w_0_300_s_0_450=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_0_450=8.67e-11
.param mcrdlm3l1_cf_w_0_300_s_0_450=5.18e-12
.param mcrdlm3l1_ca_w_0_300_s_0_600=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_0_600=7.38e-11
.param mcrdlm3l1_cf_w_0_300_s_0_600=6.84e-12
.param mcrdlm3l1_ca_w_0_300_s_0_800=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_0_800=6.09e-11
.param mcrdlm3l1_cf_w_0_300_s_0_800=8.86e-12
.param mcrdlm3l1_ca_w_0_300_s_1_000=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_1_000=5.13e-11
.param mcrdlm3l1_cf_w_0_300_s_1_000=1.09e-11
.param mcrdlm3l1_ca_w_0_300_s_1_200=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_1_200=4.41e-11
.param mcrdlm3l1_cf_w_0_300_s_1_200=1.28e-11
.param mcrdlm3l1_ca_w_0_300_s_2_100=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_2_100=2.59e-11
.param mcrdlm3l1_cf_w_0_300_s_2_100=2.04e-11
.param mcrdlm3l1_ca_w_0_300_s_3_300=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_3_300=1.51e-11
.param mcrdlm3l1_cf_w_0_300_s_3_300=2.70e-11
.param mcrdlm3l1_ca_w_0_300_s_9_000=2.37e-05
.param mcrdlm3l1_cc_w_0_300_s_9_000=2.07e-12
.param mcrdlm3l1_cf_w_0_300_s_9_000=3.80e-11
.param mcrdlm3l1_ca_w_2_400_s_0_300=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_0_300=1.23e-10
.param mcrdlm3l1_cf_w_2_400_s_0_300=3.52e-12
.param mcrdlm3l1_ca_w_2_400_s_0_360=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_0_360=1.14e-10
.param mcrdlm3l1_cf_w_2_400_s_0_360=4.20e-12
.param mcrdlm3l1_ca_w_2_400_s_0_450=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_0_450=1.03e-10
.param mcrdlm3l1_cf_w_2_400_s_0_450=5.20e-12
.param mcrdlm3l1_ca_w_2_400_s_0_600=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_0_600=8.82e-11
.param mcrdlm3l1_cf_w_2_400_s_0_600=6.83e-12
.param mcrdlm3l1_ca_w_2_400_s_0_800=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_0_800=7.31e-11
.param mcrdlm3l1_cf_w_2_400_s_0_800=8.94e-12
.param mcrdlm3l1_ca_w_2_400_s_1_000=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_1_000=6.22e-11
.param mcrdlm3l1_cf_w_2_400_s_1_000=1.10e-11
.param mcrdlm3l1_ca_w_2_400_s_1_200=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_1_200=5.38e-11
.param mcrdlm3l1_cf_w_2_400_s_1_200=1.29e-11
.param mcrdlm3l1_ca_w_2_400_s_2_100=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_2_100=3.28e-11
.param mcrdlm3l1_cf_w_2_400_s_2_100=2.05e-11
.param mcrdlm3l1_ca_w_2_400_s_3_300=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_3_300=1.97e-11
.param mcrdlm3l1_cf_w_2_400_s_3_300=2.80e-11
.param mcrdlm3l1_ca_w_2_400_s_9_000=2.37e-05
.param mcrdlm3l1_cc_w_2_400_s_9_000=3.00e-12
.param mcrdlm3l1_cf_w_2_400_s_9_000=4.15e-11
.param mcrdlm3m1_ca_w_0_300_s_0_300=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_0_300=1.01e-10
.param mcrdlm3m1_cf_w_0_300_s_0_300=5.24e-12
.param mcrdlm3m1_ca_w_0_300_s_0_360=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_0_360=9.37e-11
.param mcrdlm3m1_cf_w_0_300_s_0_360=6.25e-12
.param mcrdlm3m1_ca_w_0_300_s_0_450=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_0_450=8.35e-11
.param mcrdlm3m1_cf_w_0_300_s_0_450=7.74e-12
.param mcrdlm3m1_ca_w_0_300_s_0_600=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_0_600=7.01e-11
.param mcrdlm3m1_cf_w_0_300_s_0_600=1.01e-11
.param mcrdlm3m1_ca_w_0_300_s_0_800=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_0_800=5.70e-11
.param mcrdlm3m1_cf_w_0_300_s_0_800=1.30e-11
.param mcrdlm3m1_ca_w_0_300_s_1_000=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_1_000=4.73e-11
.param mcrdlm3m1_cf_w_0_300_s_1_000=1.58e-11
.param mcrdlm3m1_ca_w_0_300_s_1_200=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_1_200=4.00e-11
.param mcrdlm3m1_cf_w_0_300_s_1_200=1.83e-11
.param mcrdlm3m1_ca_w_0_300_s_2_100=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_2_100=2.17e-11
.param mcrdlm3m1_cf_w_0_300_s_2_100=2.77e-11
.param mcrdlm3m1_ca_w_0_300_s_3_300=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_3_300=1.18e-11
.param mcrdlm3m1_cf_w_0_300_s_3_300=3.49e-11
.param mcrdlm3m1_ca_w_0_300_s_9_000=3.64e-05
.param mcrdlm3m1_cc_w_0_300_s_9_000=1.31e-12
.param mcrdlm3m1_cf_w_0_300_s_9_000=4.43e-11
.param mcrdlm3m1_ca_w_2_400_s_0_300=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_0_300=1.17e-10
.param mcrdlm3m1_cf_w_2_400_s_0_300=5.26e-12
.param mcrdlm3m1_ca_w_2_400_s_0_360=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_0_360=1.09e-10
.param mcrdlm3m1_cf_w_2_400_s_0_360=6.27e-12
.param mcrdlm3m1_ca_w_2_400_s_0_450=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_0_450=9.80e-11
.param mcrdlm3m1_cf_w_2_400_s_0_450=7.74e-12
.param mcrdlm3m1_ca_w_2_400_s_0_600=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_0_600=8.29e-11
.param mcrdlm3m1_cf_w_2_400_s_0_600=1.01e-11
.param mcrdlm3m1_ca_w_2_400_s_0_800=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_0_800=6.80e-11
.param mcrdlm3m1_cf_w_2_400_s_0_800=1.31e-11
.param mcrdlm3m1_ca_w_2_400_s_1_000=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_1_000=5.70e-11
.param mcrdlm3m1_cf_w_2_400_s_1_000=1.59e-11
.param mcrdlm3m1_ca_w_2_400_s_1_200=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_1_200=4.88e-11
.param mcrdlm3m1_cf_w_2_400_s_1_200=1.85e-11
.param mcrdlm3m1_ca_w_2_400_s_2_100=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_2_100=2.82e-11
.param mcrdlm3m1_cf_w_2_400_s_2_100=2.79e-11
.param mcrdlm3m1_ca_w_2_400_s_3_300=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_3_300=1.61e-11
.param mcrdlm3m1_cf_w_2_400_s_3_300=3.61e-11
.param mcrdlm3m1_ca_w_2_400_s_9_000=3.64e-05
.param mcrdlm3m1_cc_w_2_400_s_9_000=2.13e-12
.param mcrdlm3m1_cf_w_2_400_s_9_000=4.82e-11
.param mcrdlm3m2_ca_w_0_300_s_0_300=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_0_300=9.31e-11
.param mcrdlm3m2_cf_w_0_300_s_0_300=1.16e-11
.param mcrdlm3m2_ca_w_0_300_s_0_360=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_0_360=8.55e-11
.param mcrdlm3m2_cf_w_0_300_s_0_360=1.36e-11
.param mcrdlm3m2_ca_w_0_300_s_0_450=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_0_450=7.53e-11
.param mcrdlm3m2_cf_w_0_300_s_0_450=1.65e-11
.param mcrdlm3m2_ca_w_0_300_s_0_600=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_0_600=6.18e-11
.param mcrdlm3m2_cf_w_0_300_s_0_600=2.09e-11
.param mcrdlm3m2_ca_w_0_300_s_0_800=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_0_800=4.88e-11
.param mcrdlm3m2_cf_w_0_300_s_0_800=2.59e-11
.param mcrdlm3m2_ca_w_0_300_s_1_000=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_1_000=3.92e-11
.param mcrdlm3m2_cf_w_0_300_s_1_000=3.02e-11
.param mcrdlm3m2_ca_w_0_300_s_1_200=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_1_200=3.23e-11
.param mcrdlm3m2_cf_w_0_300_s_1_200=3.38e-11
.param mcrdlm3m2_ca_w_0_300_s_2_100=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_2_100=1.55e-11
.param mcrdlm3m2_cf_w_0_300_s_2_100=4.52e-11
.param mcrdlm3m2_ca_w_0_300_s_3_300=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_3_300=7.64e-12
.param mcrdlm3m2_cf_w_0_300_s_3_300=5.18e-11
.param mcrdlm3m2_ca_w_0_300_s_9_000=8.57e-05
.param mcrdlm3m2_cc_w_0_300_s_9_000=7.65e-13
.param mcrdlm3m2_cf_w_0_300_s_9_000=5.84e-11
.param mcrdlm3m2_ca_w_2_400_s_0_300=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_0_300=1.07e-10
.param mcrdlm3m2_cf_w_2_400_s_0_300=1.16e-11
.param mcrdlm3m2_ca_w_2_400_s_0_360=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_0_360=9.93e-11
.param mcrdlm3m2_cf_w_2_400_s_0_360=1.37e-11
.param mcrdlm3m2_ca_w_2_400_s_0_450=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_0_450=8.82e-11
.param mcrdlm3m2_cf_w_2_400_s_0_450=1.65e-11
.param mcrdlm3m2_ca_w_2_400_s_0_600=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_0_600=7.34e-11
.param mcrdlm3m2_cf_w_2_400_s_0_600=2.09e-11
.param mcrdlm3m2_ca_w_2_400_s_0_800=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_0_800=5.89e-11
.param mcrdlm3m2_cf_w_2_400_s_0_800=2.59e-11
.param mcrdlm3m2_ca_w_2_400_s_1_000=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_1_000=4.84e-11
.param mcrdlm3m2_cf_w_2_400_s_1_000=3.03e-11
.param mcrdlm3m2_ca_w_2_400_s_1_200=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_1_200=4.05e-11
.param mcrdlm3m2_cf_w_2_400_s_1_200=3.39e-11
.param mcrdlm3m2_ca_w_2_400_s_2_100=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_2_100=2.19e-11
.param mcrdlm3m2_cf_w_2_400_s_2_100=4.54e-11
.param mcrdlm3m2_ca_w_2_400_s_3_300=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_3_300=1.18e-11
.param mcrdlm3m2_cf_w_2_400_s_3_300=5.36e-11
.param mcrdlm3m2_ca_w_2_400_s_9_000=8.57e-05
.param mcrdlm3m2_cc_w_2_400_s_9_000=1.27e-12
.param mcrdlm3m2_cf_w_2_400_s_9_000=6.34e-11
.param mcm5m4f_ca_w_0_300_s_0_300=7.70e-05
.param mcm5m4f_cc_w_0_300_s_0_300=9.38e-11
.param mcm5m4f_cf_w_0_300_s_0_300=1.01e-11
.param mcm5m4f_ca_w_0_300_s_0_360=7.70e-05
.param mcm5m4f_cc_w_0_300_s_0_360=8.64e-11
.param mcm5m4f_cf_w_0_300_s_0_360=1.20e-11
.param mcm5m4f_ca_w_0_300_s_0_450=7.70e-05
.param mcm5m4f_cc_w_0_300_s_0_450=7.58e-11
.param mcm5m4f_cf_w_0_300_s_0_450=1.47e-11
.param mcm5m4f_ca_w_0_300_s_0_600=7.70e-05
.param mcm5m4f_cc_w_0_300_s_0_600=6.20e-11
.param mcm5m4f_cf_w_0_300_s_0_600=1.88e-11
.param mcm5m4f_ca_w_0_300_s_0_800=7.70e-05
.param mcm5m4f_cc_w_0_300_s_0_800=4.84e-11
.param mcm5m4f_cf_w_0_300_s_0_800=2.37e-11
.param mcm5m4f_ca_w_0_300_s_1_000=7.70e-05
.param mcm5m4f_cc_w_0_300_s_1_000=3.85e-11
.param mcm5m4f_cf_w_0_300_s_1_000=2.80e-11
.param mcm5m4f_ca_w_0_300_s_1_200=7.70e-05
.param mcm5m4f_cc_w_0_300_s_1_200=3.12e-11
.param mcm5m4f_cf_w_0_300_s_1_200=3.17e-11
.param mcm5m4f_ca_w_0_300_s_2_100=7.70e-05
.param mcm5m4f_cc_w_0_300_s_2_100=1.39e-11
.param mcm5m4f_cf_w_0_300_s_2_100=4.31e-11
.param mcm5m4f_ca_w_0_300_s_3_300=7.70e-05
.param mcm5m4f_cc_w_0_300_s_3_300=5.70e-12
.param mcm5m4f_cf_w_0_300_s_3_300=5.01e-11
.param mcm5m4f_ca_w_0_300_s_9_000=7.70e-05
.param mcm5m4f_cc_w_0_300_s_9_000=2.30e-13
.param mcm5m4f_cf_w_0_300_s_9_000=5.53e-11
.param mcm5m4f_ca_w_2_400_s_0_300=7.70e-05
.param mcm5m4f_cc_w_2_400_s_0_300=1.04e-10
.param mcm5m4f_cf_w_2_400_s_0_300=1.02e-11
.param mcm5m4f_ca_w_2_400_s_0_360=7.70e-05
.param mcm5m4f_cc_w_2_400_s_0_360=9.57e-11
.param mcm5m4f_cf_w_2_400_s_0_360=1.21e-11
.param mcm5m4f_ca_w_2_400_s_0_450=7.70e-05
.param mcm5m4f_cc_w_2_400_s_0_450=8.47e-11
.param mcm5m4f_cf_w_2_400_s_0_450=1.47e-11
.param mcm5m4f_ca_w_2_400_s_0_600=7.70e-05
.param mcm5m4f_cc_w_2_400_s_0_600=6.97e-11
.param mcm5m4f_cf_w_2_400_s_0_600=1.89e-11
.param mcm5m4f_ca_w_2_400_s_0_800=7.70e-05
.param mcm5m4f_cc_w_2_400_s_0_800=5.49e-11
.param mcm5m4f_cf_w_2_400_s_0_800=2.38e-11
.param mcm5m4f_ca_w_2_400_s_1_000=7.70e-05
.param mcm5m4f_cc_w_2_400_s_1_000=4.39e-11
.param mcm5m4f_cf_w_2_400_s_1_000=2.81e-11
.param mcm5m4f_ca_w_2_400_s_1_200=7.70e-05
.param mcm5m4f_cc_w_2_400_s_1_200=3.59e-11
.param mcm5m4f_cf_w_2_400_s_1_200=3.19e-11
.param mcm5m4f_ca_w_2_400_s_2_100=7.70e-05
.param mcm5m4f_cc_w_2_400_s_2_100=1.70e-11
.param mcm5m4f_cf_w_2_400_s_2_100=4.38e-11
.param mcm5m4f_ca_w_2_400_s_3_300=7.70e-05
.param mcm5m4f_cc_w_2_400_s_3_300=7.38e-12
.param mcm5m4f_cf_w_2_400_s_3_300=5.17e-11
.param mcm5m4f_ca_w_2_400_s_9_000=7.70e-05
.param mcm5m4f_cc_w_2_400_s_9_000=3.05e-13
.param mcm5m4f_cf_w_2_400_s_9_000=5.85e-11
.param mcm5m4d_ca_w_0_300_s_0_300=7.78e-05
.param mcm5m4d_cc_w_0_300_s_0_300=9.36e-11
.param mcm5m4d_cf_w_0_300_s_0_300=1.02e-11
.param mcm5m4d_ca_w_0_300_s_0_360=7.78e-05
.param mcm5m4d_cc_w_0_300_s_0_360=8.61e-11
.param mcm5m4d_cf_w_0_300_s_0_360=1.21e-11
.param mcm5m4d_ca_w_0_300_s_0_450=7.78e-05
.param mcm5m4d_cc_w_0_300_s_0_450=7.56e-11
.param mcm5m4d_cf_w_0_300_s_0_450=1.48e-11
.param mcm5m4d_ca_w_0_300_s_0_600=7.78e-05
.param mcm5m4d_cc_w_0_300_s_0_600=6.17e-11
.param mcm5m4d_cf_w_0_300_s_0_600=1.90e-11
.param mcm5m4d_ca_w_0_300_s_0_800=7.78e-05
.param mcm5m4d_cc_w_0_300_s_0_800=4.82e-11
.param mcm5m4d_cf_w_0_300_s_0_800=2.39e-11
.param mcm5m4d_ca_w_0_300_s_1_000=7.78e-05
.param mcm5m4d_cc_w_0_300_s_1_000=3.82e-11
.param mcm5m4d_cf_w_0_300_s_1_000=2.83e-11
.param mcm5m4d_ca_w_0_300_s_1_200=7.78e-05
.param mcm5m4d_cc_w_0_300_s_1_200=3.08e-11
.param mcm5m4d_cf_w_0_300_s_1_200=3.21e-11
.param mcm5m4d_ca_w_0_300_s_2_100=7.78e-05
.param mcm5m4d_cc_w_0_300_s_2_100=1.35e-11
.param mcm5m4d_cf_w_0_300_s_2_100=4.36e-11
.param mcm5m4d_ca_w_0_300_s_3_300=7.78e-05
.param mcm5m4d_cc_w_0_300_s_3_300=5.39e-12
.param mcm5m4d_cf_w_0_300_s_3_300=5.04e-11
.param mcm5m4d_ca_w_0_300_s_9_000=7.78e-05
.param mcm5m4d_cc_w_0_300_s_9_000=1.45e-13
.param mcm5m4d_cf_w_0_300_s_9_000=5.54e-11
.param mcm5m4d_ca_w_2_400_s_0_300=7.78e-05
.param mcm5m4d_cc_w_2_400_s_0_300=1.04e-10
.param mcm5m4d_cf_w_2_400_s_0_300=1.03e-11
.param mcm5m4d_ca_w_2_400_s_0_360=7.78e-05
.param mcm5m4d_cc_w_2_400_s_0_360=9.52e-11
.param mcm5m4d_cf_w_2_400_s_0_360=1.22e-11
.param mcm5m4d_ca_w_2_400_s_0_450=7.78e-05
.param mcm5m4d_cc_w_2_400_s_0_450=8.40e-11
.param mcm5m4d_cf_w_2_400_s_0_450=1.49e-11
.param mcm5m4d_ca_w_2_400_s_0_600=7.78e-05
.param mcm5m4d_cc_w_2_400_s_0_600=6.90e-11
.param mcm5m4d_cf_w_2_400_s_0_600=1.91e-11
.param mcm5m4d_ca_w_2_400_s_0_800=7.78e-05
.param mcm5m4d_cc_w_2_400_s_0_800=5.42e-11
.param mcm5m4d_cf_w_2_400_s_0_800=2.41e-11
.param mcm5m4d_ca_w_2_400_s_1_000=7.78e-05
.param mcm5m4d_cc_w_2_400_s_1_000=4.33e-11
.param mcm5m4d_cf_w_2_400_s_1_000=2.85e-11
.param mcm5m4d_ca_w_2_400_s_1_200=7.78e-05
.param mcm5m4d_cc_w_2_400_s_1_200=3.52e-11
.param mcm5m4d_cf_w_2_400_s_1_200=3.23e-11
.param mcm5m4d_ca_w_2_400_s_2_100=7.78e-05
.param mcm5m4d_cc_w_2_400_s_2_100=1.63e-11
.param mcm5m4d_cf_w_2_400_s_2_100=4.42e-11
.param mcm5m4d_ca_w_2_400_s_3_300=7.78e-05
.param mcm5m4d_cc_w_2_400_s_3_300=6.86e-12
.param mcm5m4d_cf_w_2_400_s_3_300=5.20e-11
.param mcm5m4d_ca_w_2_400_s_9_000=7.78e-05
.param mcm5m4d_cc_w_2_400_s_9_000=2.25e-13
.param mcm5m4d_cf_w_2_400_s_9_000=5.84e-11
.param mcm5m4p1_ca_w_0_300_s_0_300=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_0_300=9.34e-11
.param mcm5m4p1_cf_w_0_300_s_0_300=1.03e-11
.param mcm5m4p1_ca_w_0_300_s_0_360=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_0_360=8.59e-11
.param mcm5m4p1_cf_w_0_300_s_0_360=1.22e-11
.param mcm5m4p1_ca_w_0_300_s_0_450=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_0_450=7.54e-11
.param mcm5m4p1_cf_w_0_300_s_0_450=1.50e-11
.param mcm5m4p1_ca_w_0_300_s_0_600=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_0_600=6.15e-11
.param mcm5m4p1_cf_w_0_300_s_0_600=1.92e-11
.param mcm5m4p1_ca_w_0_300_s_0_800=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_0_800=4.79e-11
.param mcm5m4p1_cf_w_0_300_s_0_800=2.42e-11
.param mcm5m4p1_ca_w_0_300_s_1_000=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_1_000=3.78e-11
.param mcm5m4p1_cf_w_0_300_s_1_000=2.86e-11
.param mcm5m4p1_ca_w_0_300_s_1_200=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_1_200=3.04e-11
.param mcm5m4p1_cf_w_0_300_s_1_200=3.24e-11
.param mcm5m4p1_ca_w_0_300_s_2_100=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_2_100=1.32e-11
.param mcm5m4p1_cf_w_0_300_s_2_100=4.40e-11
.param mcm5m4p1_ca_w_0_300_s_3_300=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_3_300=5.10e-12
.param mcm5m4p1_cf_w_0_300_s_3_300=5.08e-11
.param mcm5m4p1_ca_w_0_300_s_9_000=7.85e-05
.param mcm5m4p1_cc_w_0_300_s_9_000=1.45e-13
.param mcm5m4p1_cf_w_0_300_s_9_000=5.56e-11
.param mcm5m4p1_ca_w_2_400_s_0_300=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_0_300=1.03e-10
.param mcm5m4p1_cf_w_2_400_s_0_300=1.04e-11
.param mcm5m4p1_ca_w_2_400_s_0_360=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_0_360=9.46e-11
.param mcm5m4p1_cf_w_2_400_s_0_360=1.23e-11
.param mcm5m4p1_ca_w_2_400_s_0_450=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_0_450=8.33e-11
.param mcm5m4p1_cf_w_2_400_s_0_450=1.50e-11
.param mcm5m4p1_ca_w_2_400_s_0_600=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_0_600=6.83e-11
.param mcm5m4p1_cf_w_2_400_s_0_600=1.93e-11
.param mcm5m4p1_ca_w_2_400_s_0_800=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_0_800=5.35e-11
.param mcm5m4p1_cf_w_2_400_s_0_800=2.44e-11
.param mcm5m4p1_ca_w_2_400_s_1_000=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_1_000=4.26e-11
.param mcm5m4p1_cf_w_2_400_s_1_000=2.88e-11
.param mcm5m4p1_ca_w_2_400_s_1_200=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_1_200=3.45e-11
.param mcm5m4p1_cf_w_2_400_s_1_200=3.26e-11
.param mcm5m4p1_ca_w_2_400_s_2_100=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_2_100=1.57e-11
.param mcm5m4p1_cf_w_2_400_s_2_100=4.47e-11
.param mcm5m4p1_ca_w_2_400_s_3_300=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_3_300=6.43e-12
.param mcm5m4p1_cf_w_2_400_s_3_300=5.24e-11
.param mcm5m4p1_ca_w_2_400_s_9_000=7.85e-05
.param mcm5m4p1_cc_w_2_400_s_9_000=1.70e-13
.param mcm5m4p1_cf_w_2_400_s_9_000=5.84e-11
.param mcm5m4l1_ca_w_0_300_s_0_300=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_0_300=9.30e-11
.param mcm5m4l1_cf_w_0_300_s_0_300=1.05e-11
.param mcm5m4l1_ca_w_0_300_s_0_360=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_0_360=8.55e-11
.param mcm5m4l1_cf_w_0_300_s_0_360=1.25e-11
.param mcm5m4l1_ca_w_0_300_s_0_450=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_0_450=7.50e-11
.param mcm5m4l1_cf_w_0_300_s_0_450=1.53e-11
.param mcm5m4l1_ca_w_0_300_s_0_600=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_0_600=6.08e-11
.param mcm5m4l1_cf_w_0_300_s_0_600=1.97e-11
.param mcm5m4l1_ca_w_0_300_s_0_800=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_0_800=4.72e-11
.param mcm5m4l1_cf_w_0_300_s_0_800=2.48e-11
.param mcm5m4l1_ca_w_0_300_s_1_000=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_1_000=3.71e-11
.param mcm5m4l1_cf_w_0_300_s_1_000=2.92e-11
.param mcm5m4l1_ca_w_0_300_s_1_200=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_1_200=2.96e-11
.param mcm5m4l1_cf_w_0_300_s_1_200=3.31e-11
.param mcm5m4l1_ca_w_0_300_s_2_100=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_2_100=1.24e-11
.param mcm5m4l1_cf_w_0_300_s_2_100=4.48e-11
.param mcm5m4l1_ca_w_0_300_s_3_300=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_3_300=4.60e-12
.param mcm5m4l1_cf_w_0_300_s_3_300=5.15e-11
.param mcm5m4l1_ca_w_0_300_s_9_000=8.01e-05
.param mcm5m4l1_cc_w_0_300_s_9_000=1.60e-13
.param mcm5m4l1_cf_w_0_300_s_9_000=5.59e-11
.param mcm5m4l1_ca_w_2_400_s_0_300=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_0_300=1.02e-10
.param mcm5m4l1_cf_w_2_400_s_0_300=1.06e-11
.param mcm5m4l1_ca_w_2_400_s_0_360=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_0_360=9.33e-11
.param mcm5m4l1_cf_w_2_400_s_0_360=1.26e-11
.param mcm5m4l1_ca_w_2_400_s_0_450=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_0_450=8.20e-11
.param mcm5m4l1_cf_w_2_400_s_0_450=1.54e-11
.param mcm5m4l1_ca_w_2_400_s_0_600=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_0_600=6.70e-11
.param mcm5m4l1_cf_w_2_400_s_0_600=1.97e-11
.param mcm5m4l1_ca_w_2_400_s_0_800=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_0_800=5.22e-11
.param mcm5m4l1_cf_w_2_400_s_0_800=2.49e-11
.param mcm5m4l1_ca_w_2_400_s_1_000=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_1_000=4.12e-11
.param mcm5m4l1_cf_w_2_400_s_1_000=2.95e-11
.param mcm5m4l1_ca_w_2_400_s_1_200=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_1_200=3.32e-11
.param mcm5m4l1_cf_w_2_400_s_1_200=3.34e-11
.param mcm5m4l1_ca_w_2_400_s_2_100=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_2_100=1.45e-11
.param mcm5m4l1_cf_w_2_400_s_2_100=4.56e-11
.param mcm5m4l1_ca_w_2_400_s_3_300=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_3_300=5.55e-12
.param mcm5m4l1_cf_w_2_400_s_3_300=5.31e-11
.param mcm5m4l1_ca_w_2_400_s_9_000=8.01e-05
.param mcm5m4l1_cc_w_2_400_s_9_000=8.50e-14
.param mcm5m4l1_cf_w_2_400_s_9_000=5.84e-11
.param mcm5m4m1_ca_w_0_300_s_0_300=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_0_300=9.22e-11
.param mcm5m4m1_cf_w_0_300_s_0_300=1.10e-11
.param mcm5m4m1_ca_w_0_300_s_0_360=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_0_360=8.45e-11
.param mcm5m4m1_cf_w_0_300_s_0_360=1.31e-11
.param mcm5m4m1_ca_w_0_300_s_0_450=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_0_450=7.40e-11
.param mcm5m4m1_cf_w_0_300_s_0_450=1.60e-11
.param mcm5m4m1_ca_w_0_300_s_0_600=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_0_600=5.97e-11
.param mcm5m4m1_cf_w_0_300_s_0_600=2.06e-11
.param mcm5m4m1_ca_w_0_300_s_0_800=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_0_800=4.59e-11
.param mcm5m4m1_cf_w_0_300_s_0_800=2.60e-11
.param mcm5m4m1_ca_w_0_300_s_1_000=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_1_000=3.56e-11
.param mcm5m4m1_cf_w_0_300_s_1_000=3.07e-11
.param mcm5m4m1_ca_w_0_300_s_1_200=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_1_200=2.81e-11
.param mcm5m4m1_cf_w_0_300_s_1_200=3.48e-11
.param mcm5m4m1_ca_w_0_300_s_2_100=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_2_100=1.10e-11
.param mcm5m4m1_cf_w_0_300_s_2_100=4.66e-11
.param mcm5m4m1_ca_w_0_300_s_3_300=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_3_300=3.61e-12
.param mcm5m4m1_cf_w_0_300_s_3_300=5.31e-11
.param mcm5m4m1_ca_w_0_300_s_9_000=8.35e-05
.param mcm5m4m1_cc_w_0_300_s_9_000=5.50e-14
.param mcm5m4m1_cf_w_0_300_s_9_000=5.67e-11
.param mcm5m4m1_ca_w_2_400_s_0_300=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_0_300=9.94e-11
.param mcm5m4m1_cf_w_2_400_s_0_300=1.11e-11
.param mcm5m4m1_ca_w_2_400_s_0_360=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_0_360=9.08e-11
.param mcm5m4m1_cf_w_2_400_s_0_360=1.31e-11
.param mcm5m4m1_ca_w_2_400_s_0_450=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_0_450=7.95e-11
.param mcm5m4m1_cf_w_2_400_s_0_450=1.61e-11
.param mcm5m4m1_ca_w_2_400_s_0_600=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_0_600=6.45e-11
.param mcm5m4m1_cf_w_2_400_s_0_600=2.07e-11
.param mcm5m4m1_ca_w_2_400_s_0_800=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_0_800=4.96e-11
.param mcm5m4m1_cf_w_2_400_s_0_800=2.61e-11
.param mcm5m4m1_ca_w_2_400_s_1_000=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_1_000=3.87e-11
.param mcm5m4m1_cf_w_2_400_s_1_000=3.09e-11
.param mcm5m4m1_ca_w_2_400_s_1_200=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_1_200=3.07e-11
.param mcm5m4m1_cf_w_2_400_s_1_200=3.50e-11
.param mcm5m4m1_ca_w_2_400_s_2_100=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_2_100=1.23e-11
.param mcm5m4m1_cf_w_2_400_s_2_100=4.74e-11
.param mcm5m4m1_ca_w_2_400_s_3_300=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_3_300=4.21e-12
.param mcm5m4m1_cf_w_2_400_s_3_300=5.45e-11
.param mcm5m4m1_ca_w_2_400_s_9_000=8.35e-05
.param mcm5m4m1_cc_w_2_400_s_9_000=9.50e-14
.param mcm5m4m1_cf_w_2_400_s_9_000=5.86e-11
.param mcm5m4m2_ca_w_0_300_s_0_300=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_0_300=9.10e-11
.param mcm5m4m2_cf_w_0_300_s_0_300=1.19e-11
.param mcm5m4m2_ca_w_0_300_s_0_360=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_0_360=8.30e-11
.param mcm5m4m2_cf_w_0_300_s_0_360=1.41e-11
.param mcm5m4m2_ca_w_0_300_s_0_450=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_0_450=7.24e-11
.param mcm5m4m2_cf_w_0_300_s_0_450=1.73e-11
.param mcm5m4m2_ca_w_0_300_s_0_600=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_0_600=5.78e-11
.param mcm5m4m2_cf_w_0_300_s_0_600=2.22e-11
.param mcm5m4m2_ca_w_0_300_s_0_800=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_0_800=4.38e-11
.param mcm5m4m2_cf_w_0_300_s_0_800=2.79e-11
.param mcm5m4m2_ca_w_0_300_s_1_000=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_1_000=3.35e-11
.param mcm5m4m2_cf_w_0_300_s_1_000=3.30e-11
.param mcm5m4m2_ca_w_0_300_s_1_200=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_1_200=2.59e-11
.param mcm5m4m2_cf_w_0_300_s_1_200=3.73e-11
.param mcm5m4m2_ca_w_0_300_s_2_100=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_2_100=9.12e-12
.param mcm5m4m2_cf_w_0_300_s_2_100=4.94e-11
.param mcm5m4m2_ca_w_0_300_s_3_300=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_3_300=2.55e-12
.param mcm5m4m2_cf_w_0_300_s_3_300=5.55e-11
.param mcm5m4m2_ca_w_0_300_s_9_000=8.92e-05
.param mcm5m4m2_cc_w_0_300_s_9_000=4.00e-14
.param mcm5m4m2_cf_w_0_300_s_9_000=5.80e-11
.param mcm5m4m2_ca_w_2_400_s_0_300=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_0_300=9.61e-11
.param mcm5m4m2_cf_w_2_400_s_0_300=1.19e-11
.param mcm5m4m2_ca_w_2_400_s_0_360=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_0_360=8.77e-11
.param mcm5m4m2_cf_w_2_400_s_0_360=1.41e-11
.param mcm5m4m2_ca_w_2_400_s_0_450=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_0_450=7.62e-11
.param mcm5m4m2_cf_w_2_400_s_0_450=1.73e-11
.param mcm5m4m2_ca_w_2_400_s_0_600=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_0_600=6.12e-11
.param mcm5m4m2_cf_w_2_400_s_0_600=2.22e-11
.param mcm5m4m2_ca_w_2_400_s_0_800=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_0_800=4.63e-11
.param mcm5m4m2_cf_w_2_400_s_0_800=2.81e-11
.param mcm5m4m2_ca_w_2_400_s_1_000=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_1_000=3.54e-11
.param mcm5m4m2_cf_w_2_400_s_1_000=3.32e-11
.param mcm5m4m2_ca_w_2_400_s_1_200=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_1_200=2.75e-11
.param mcm5m4m2_cf_w_2_400_s_1_200=3.76e-11
.param mcm5m4m2_ca_w_2_400_s_2_100=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_2_100=9.85e-12
.param mcm5m4m2_cf_w_2_400_s_2_100=5.03e-11
.param mcm5m4m2_ca_w_2_400_s_3_300=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_3_300=2.76e-12
.param mcm5m4m2_cf_w_2_400_s_3_300=5.66e-11
.param mcm5m4m2_ca_w_2_400_s_9_000=8.92e-05
.param mcm5m4m2_cc_w_2_400_s_9_000=5.00e-15
.param mcm5m4m2_cf_w_2_400_s_9_000=5.94e-11
.param mcm5m4m3_ca_w_0_300_s_0_300=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_0_300=7.96e-11
.param mcm5m4m3_cf_w_0_300_s_0_300=2.07e-11
.param mcm5m4m3_ca_w_0_300_s_0_360=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_0_360=7.11e-11
.param mcm5m4m3_cf_w_0_300_s_0_360=2.43e-11
.param mcm5m4m3_ca_w_0_300_s_0_450=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_0_450=6.04e-11
.param mcm5m4m3_cf_w_0_300_s_0_450=2.95e-11
.param mcm5m4m3_ca_w_0_300_s_0_600=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_0_600=4.57e-11
.param mcm5m4m3_cf_w_0_300_s_0_600=3.72e-11
.param mcm5m4m3_ca_w_0_300_s_0_800=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_0_800=3.16e-11
.param mcm5m4m3_cf_w_0_300_s_0_800=4.58e-11
.param mcm5m4m3_ca_w_0_300_s_1_000=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_1_000=2.17e-11
.param mcm5m4m3_cf_w_0_300_s_1_000=5.29e-11
.param mcm5m4m3_ca_w_0_300_s_1_200=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_1_200=1.49e-11
.param mcm5m4m3_cf_w_0_300_s_1_200=5.81e-11
.param mcm5m4m3_ca_w_0_300_s_2_100=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_2_100=2.94e-12
.param mcm5m4m3_cf_w_0_300_s_2_100=6.87e-11
.param mcm5m4m3_ca_w_0_300_s_3_300=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_3_300=4.25e-13
.param mcm5m4m3_cf_w_0_300_s_3_300=7.12e-11
.param mcm5m4m3_ca_w_0_300_s_9_000=1.57e-04
.param mcm5m4m3_cc_w_0_300_s_9_000=0.00e+00
.param mcm5m4m3_cf_w_0_300_s_9_000=7.16e-11
.param mcm5m4m3_ca_w_2_400_s_0_300=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_0_300=8.05e-11
.param mcm5m4m3_cf_w_2_400_s_0_300=2.07e-11
.param mcm5m4m3_ca_w_2_400_s_0_360=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_0_360=7.21e-11
.param mcm5m4m3_cf_w_2_400_s_0_360=2.44e-11
.param mcm5m4m3_ca_w_2_400_s_0_450=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_0_450=6.07e-11
.param mcm5m4m3_cf_w_2_400_s_0_450=2.95e-11
.param mcm5m4m3_ca_w_2_400_s_0_600=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_0_600=4.63e-11
.param mcm5m4m3_cf_w_2_400_s_0_600=3.72e-11
.param mcm5m4m3_ca_w_2_400_s_0_800=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_0_800=3.18e-11
.param mcm5m4m3_cf_w_2_400_s_0_800=4.60e-11
.param mcm5m4m3_ca_w_2_400_s_1_000=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_1_000=2.19e-11
.param mcm5m4m3_cf_w_2_400_s_1_000=5.28e-11
.param mcm5m4m3_ca_w_2_400_s_1_200=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_1_200=1.50e-11
.param mcm5m4m3_cf_w_2_400_s_1_200=5.81e-11
.param mcm5m4m3_ca_w_2_400_s_2_100=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_2_100=2.95e-12
.param mcm5m4m3_cf_w_2_400_s_2_100=6.90e-11
.param mcm5m4m3_ca_w_2_400_s_3_300=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_3_300=4.00e-13
.param mcm5m4m3_cf_w_2_400_s_3_300=7.16e-11
.param mcm5m4m3_ca_w_2_400_s_9_000=1.57e-04
.param mcm5m4m3_cc_w_2_400_s_9_000=5.00e-14
.param mcm5m4m3_cf_w_2_400_s_9_000=7.21e-11
.param mcrdlm4f_ca_w_0_300_s_0_300=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_0_300=1.07e-10
.param mcrdlm4f_cf_w_0_300_s_0_300=1.88e-12
.param mcrdlm4f_ca_w_0_300_s_0_360=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_0_360=1.00e-10
.param mcrdlm4f_cf_w_0_300_s_0_360=2.25e-12
.param mcrdlm4f_ca_w_0_300_s_0_450=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_0_450=9.09e-11
.param mcrdlm4f_cf_w_0_300_s_0_450=2.84e-12
.param mcrdlm4f_ca_w_0_300_s_0_600=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_0_600=7.80e-11
.param mcrdlm4f_cf_w_0_300_s_0_600=3.80e-12
.param mcrdlm4f_ca_w_0_300_s_0_800=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_0_800=6.61e-11
.param mcrdlm4f_cf_w_0_300_s_0_800=4.91e-12
.param mcrdlm4f_ca_w_0_300_s_1_000=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_1_000=5.70e-11
.param mcrdlm4f_cf_w_0_300_s_1_000=6.09e-12
.param mcrdlm4f_ca_w_0_300_s_1_200=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_1_200=5.01e-11
.param mcrdlm4f_cf_w_0_300_s_1_200=7.24e-12
.param mcrdlm4f_ca_w_0_300_s_2_100=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_2_100=3.25e-11
.param mcrdlm4f_cf_w_0_300_s_2_100=1.22e-11
.param mcrdlm4f_ca_w_0_300_s_3_300=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_3_300=2.13e-11
.param mcrdlm4f_cf_w_0_300_s_3_300=1.72e-11
.param mcrdlm4f_ca_w_0_300_s_9_000=1.27e-05
.param mcrdlm4f_cc_w_0_300_s_9_000=4.11e-12
.param mcrdlm4f_cf_w_0_300_s_9_000=2.94e-11
.param mcrdlm4f_ca_w_2_400_s_0_300=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_0_300=1.32e-10
.param mcrdlm4f_cf_w_2_400_s_0_300=1.90e-12
.param mcrdlm4f_ca_w_2_400_s_0_360=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_0_360=1.24e-10
.param mcrdlm4f_cf_w_2_400_s_0_360=2.28e-12
.param mcrdlm4f_ca_w_2_400_s_0_450=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_0_450=1.13e-10
.param mcrdlm4f_cf_w_2_400_s_0_450=2.83e-12
.param mcrdlm4f_ca_w_2_400_s_0_600=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_0_600=9.74e-11
.param mcrdlm4f_cf_w_2_400_s_0_600=3.75e-12
.param mcrdlm4f_ca_w_2_400_s_0_800=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_0_800=8.23e-11
.param mcrdlm4f_cf_w_2_400_s_0_800=4.96e-12
.param mcrdlm4f_ca_w_2_400_s_1_000=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_1_000=7.12e-11
.param mcrdlm4f_cf_w_2_400_s_1_000=6.14e-12
.param mcrdlm4f_ca_w_2_400_s_1_200=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_1_200=6.27e-11
.param mcrdlm4f_cf_w_2_400_s_1_200=7.31e-12
.param mcrdlm4f_ca_w_2_400_s_2_100=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_2_100=4.09e-11
.param mcrdlm4f_cf_w_2_400_s_2_100=1.22e-11
.param mcrdlm4f_ca_w_2_400_s_3_300=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_3_300=2.67e-11
.param mcrdlm4f_cf_w_2_400_s_3_300=1.78e-11
.param mcrdlm4f_ca_w_2_400_s_9_000=1.27e-05
.param mcrdlm4f_cc_w_2_400_s_9_000=5.36e-12
.param mcrdlm4f_cf_w_2_400_s_9_000=3.22e-11
.param mcrdlm4d_ca_w_0_300_s_0_300=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_0_300=1.07e-10
.param mcrdlm4d_cf_w_0_300_s_0_300=1.98e-12
.param mcrdlm4d_ca_w_0_300_s_0_360=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_0_360=9.98e-11
.param mcrdlm4d_cf_w_0_300_s_0_360=2.38e-12
.param mcrdlm4d_ca_w_0_300_s_0_450=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_0_450=9.07e-11
.param mcrdlm4d_cf_w_0_300_s_0_450=3.00e-12
.param mcrdlm4d_ca_w_0_300_s_0_600=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_0_600=7.78e-11
.param mcrdlm4d_cf_w_0_300_s_0_600=4.02e-12
.param mcrdlm4d_ca_w_0_300_s_0_800=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_0_800=6.58e-11
.param mcrdlm4d_cf_w_0_300_s_0_800=5.19e-12
.param mcrdlm4d_ca_w_0_300_s_1_000=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_1_000=5.66e-11
.param mcrdlm4d_cf_w_0_300_s_1_000=6.42e-12
.param mcrdlm4d_ca_w_0_300_s_1_200=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_1_200=4.97e-11
.param mcrdlm4d_cf_w_0_300_s_1_200=7.63e-12
.param mcrdlm4d_ca_w_0_300_s_2_100=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_2_100=3.19e-11
.param mcrdlm4d_cf_w_0_300_s_2_100=1.28e-11
.param mcrdlm4d_ca_w_0_300_s_3_300=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_3_300=2.07e-11
.param mcrdlm4d_cf_w_0_300_s_3_300=1.80e-11
.param mcrdlm4d_ca_w_0_300_s_9_000=1.34e-05
.param mcrdlm4d_cc_w_0_300_s_9_000=3.82e-12
.param mcrdlm4d_cf_w_0_300_s_9_000=3.02e-11
.param mcrdlm4d_ca_w_2_400_s_0_300=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_0_300=1.31e-10
.param mcrdlm4d_cf_w_2_400_s_0_300=2.01e-12
.param mcrdlm4d_ca_w_2_400_s_0_360=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_0_360=1.23e-10
.param mcrdlm4d_cf_w_2_400_s_0_360=2.41e-12
.param mcrdlm4d_ca_w_2_400_s_0_450=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_0_450=1.12e-10
.param mcrdlm4d_cf_w_2_400_s_0_450=3.00e-12
.param mcrdlm4d_ca_w_2_400_s_0_600=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_0_600=9.68e-11
.param mcrdlm4d_cf_w_2_400_s_0_600=3.97e-12
.param mcrdlm4d_ca_w_2_400_s_0_800=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_0_800=8.15e-11
.param mcrdlm4d_cf_w_2_400_s_0_800=5.24e-12
.param mcrdlm4d_ca_w_2_400_s_1_000=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_1_000=7.05e-11
.param mcrdlm4d_cf_w_2_400_s_1_000=6.49e-12
.param mcrdlm4d_ca_w_2_400_s_1_200=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_1_200=6.20e-11
.param mcrdlm4d_cf_w_2_400_s_1_200=7.71e-12
.param mcrdlm4d_ca_w_2_400_s_2_100=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_2_100=4.01e-11
.param mcrdlm4d_cf_w_2_400_s_2_100=1.28e-11
.param mcrdlm4d_ca_w_2_400_s_3_300=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_3_300=2.59e-11
.param mcrdlm4d_cf_w_2_400_s_3_300=1.86e-11
.param mcrdlm4d_ca_w_2_400_s_9_000=1.34e-05
.param mcrdlm4d_cc_w_2_400_s_9_000=4.98e-12
.param mcrdlm4d_cf_w_2_400_s_9_000=3.31e-11
.param mcrdlm4p1_ca_w_0_300_s_0_300=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_0_300=1.07e-10
.param mcrdlm4p1_cf_w_0_300_s_0_300=2.09e-12
.param mcrdlm4p1_ca_w_0_300_s_0_360=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_0_360=9.96e-11
.param mcrdlm4p1_cf_w_0_300_s_0_360=2.51e-12
.param mcrdlm4p1_ca_w_0_300_s_0_450=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_0_450=9.03e-11
.param mcrdlm4p1_cf_w_0_300_s_0_450=3.16e-12
.param mcrdlm4p1_ca_w_0_300_s_0_600=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_0_600=7.75e-11
.param mcrdlm4p1_cf_w_0_300_s_0_600=4.23e-12
.param mcrdlm4p1_ca_w_0_300_s_0_800=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_0_800=6.54e-11
.param mcrdlm4p1_cf_w_0_300_s_0_800=5.46e-12
.param mcrdlm4p1_ca_w_0_300_s_1_000=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_1_000=5.63e-11
.param mcrdlm4p1_cf_w_0_300_s_1_000=6.76e-12
.param mcrdlm4p1_ca_w_0_300_s_1_200=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_1_200=4.93e-11
.param mcrdlm4p1_cf_w_0_300_s_1_200=8.01e-12
.param mcrdlm4p1_ca_w_0_300_s_2_100=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_2_100=3.14e-11
.param mcrdlm4p1_cf_w_0_300_s_2_100=1.34e-11
.param mcrdlm4p1_ca_w_0_300_s_3_300=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_3_300=2.02e-11
.param mcrdlm4p1_cf_w_0_300_s_3_300=1.88e-11
.param mcrdlm4p1_ca_w_0_300_s_9_000=1.41e-05
.param mcrdlm4p1_cc_w_0_300_s_9_000=3.56e-12
.param mcrdlm4p1_cf_w_0_300_s_9_000=3.09e-11
.param mcrdlm4p1_ca_w_2_400_s_0_300=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_0_300=1.31e-10
.param mcrdlm4p1_cf_w_2_400_s_0_300=2.13e-12
.param mcrdlm4p1_ca_w_2_400_s_0_360=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_0_360=1.22e-10
.param mcrdlm4p1_cf_w_2_400_s_0_360=2.55e-12
.param mcrdlm4p1_ca_w_2_400_s_0_450=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_0_450=1.11e-10
.param mcrdlm4p1_cf_w_2_400_s_0_450=3.17e-12
.param mcrdlm4p1_ca_w_2_400_s_0_600=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_0_600=9.61e-11
.param mcrdlm4p1_cf_w_2_400_s_0_600=4.18e-12
.param mcrdlm4p1_ca_w_2_400_s_0_800=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_0_800=8.09e-11
.param mcrdlm4p1_cf_w_2_400_s_0_800=5.52e-12
.param mcrdlm4p1_ca_w_2_400_s_1_000=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_1_000=6.97e-11
.param mcrdlm4p1_cf_w_2_400_s_1_000=6.83e-12
.param mcrdlm4p1_ca_w_2_400_s_1_200=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_1_200=6.13e-11
.param mcrdlm4p1_cf_w_2_400_s_1_200=8.11e-12
.param mcrdlm4p1_ca_w_2_400_s_2_100=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_2_100=3.94e-11
.param mcrdlm4p1_cf_w_2_400_s_2_100=1.34e-11
.param mcrdlm4p1_ca_w_2_400_s_3_300=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_3_300=2.52e-11
.param mcrdlm4p1_cf_w_2_400_s_3_300=1.94e-11
.param mcrdlm4p1_ca_w_2_400_s_9_000=1.41e-05
.param mcrdlm4p1_cc_w_2_400_s_9_000=4.65e-12
.param mcrdlm4p1_cf_w_2_400_s_9_000=3.39e-11
.param mcrdlm4l1_ca_w_0_300_s_0_300=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_0_300=1.06e-10
.param mcrdlm4l1_cf_w_0_300_s_0_300=2.32e-12
.param mcrdlm4l1_ca_w_0_300_s_0_360=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_0_360=9.92e-11
.param mcrdlm4l1_cf_w_0_300_s_0_360=2.78e-12
.param mcrdlm4l1_ca_w_0_300_s_0_450=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_0_450=8.98e-11
.param mcrdlm4l1_cf_w_0_300_s_0_450=3.49e-12
.param mcrdlm4l1_ca_w_0_300_s_0_600=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_0_600=7.71e-11
.param mcrdlm4l1_cf_w_0_300_s_0_600=4.67e-12
.param mcrdlm4l1_ca_w_0_300_s_0_800=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_0_800=6.47e-11
.param mcrdlm4l1_cf_w_0_300_s_0_800=6.04e-12
.param mcrdlm4l1_ca_w_0_300_s_1_000=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_1_000=5.55e-11
.param mcrdlm4l1_cf_w_0_300_s_1_000=7.46e-12
.param mcrdlm4l1_ca_w_0_300_s_1_200=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_1_200=4.86e-11
.param mcrdlm4l1_cf_w_0_300_s_1_200=8.84e-12
.param mcrdlm4l1_ca_w_0_300_s_2_100=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_2_100=3.04e-11
.param mcrdlm4l1_cf_w_0_300_s_2_100=1.46e-11
.param mcrdlm4l1_ca_w_0_300_s_3_300=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_3_300=1.91e-11
.param mcrdlm4l1_cf_w_0_300_s_3_300=2.03e-11
.param mcrdlm4l1_ca_w_0_300_s_9_000=1.57e-05
.param mcrdlm4l1_cc_w_0_300_s_9_000=3.08e-12
.param mcrdlm4l1_cf_w_0_300_s_9_000=3.25e-11
.param mcrdlm4l1_ca_w_2_400_s_0_300=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_0_300=1.29e-10
.param mcrdlm4l1_cf_w_2_400_s_0_300=2.34e-12
.param mcrdlm4l1_ca_w_2_400_s_0_360=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_0_360=1.21e-10
.param mcrdlm4l1_cf_w_2_400_s_0_360=2.80e-12
.param mcrdlm4l1_ca_w_2_400_s_0_450=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_0_450=1.10e-10
.param mcrdlm4l1_cf_w_2_400_s_0_450=3.49e-12
.param mcrdlm4l1_ca_w_2_400_s_0_600=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_0_600=9.46e-11
.param mcrdlm4l1_cf_w_2_400_s_0_600=4.61e-12
.param mcrdlm4l1_ca_w_2_400_s_0_800=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_0_800=7.96e-11
.param mcrdlm4l1_cf_w_2_400_s_0_800=6.08e-12
.param mcrdlm4l1_ca_w_2_400_s_1_000=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_1_000=6.84e-11
.param mcrdlm4l1_cf_w_2_400_s_1_000=7.53e-12
.param mcrdlm4l1_ca_w_2_400_s_1_200=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_1_200=5.98e-11
.param mcrdlm4l1_cf_w_2_400_s_1_200=8.92e-12
.param mcrdlm4l1_ca_w_2_400_s_2_100=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_2_100=3.80e-11
.param mcrdlm4l1_cf_w_2_400_s_2_100=1.47e-11
.param mcrdlm4l1_ca_w_2_400_s_3_300=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_3_300=2.39e-11
.param mcrdlm4l1_cf_w_2_400_s_3_300=2.11e-11
.param mcrdlm4l1_ca_w_2_400_s_9_000=1.57e-05
.param mcrdlm4l1_cc_w_2_400_s_9_000=4.05e-12
.param mcrdlm4l1_cf_w_2_400_s_9_000=3.55e-11
.param mcrdlm4m1_ca_w_0_300_s_0_300=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_0_300=1.06e-10
.param mcrdlm4m1_cf_w_0_300_s_0_300=2.81e-12
.param mcrdlm4m1_ca_w_0_300_s_0_360=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_0_360=9.83e-11
.param mcrdlm4m1_cf_w_0_300_s_0_360=3.36e-12
.param mcrdlm4m1_ca_w_0_300_s_0_450=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_0_450=8.89e-11
.param mcrdlm4m1_cf_w_0_300_s_0_450=4.22e-12
.param mcrdlm4m1_ca_w_0_300_s_0_600=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_0_600=7.61e-11
.param mcrdlm4m1_cf_w_0_300_s_0_600=5.60e-12
.param mcrdlm4m1_ca_w_0_300_s_0_800=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_0_800=6.34e-11
.param mcrdlm4m1_cf_w_0_300_s_0_800=7.26e-12
.param mcrdlm4m1_ca_w_0_300_s_1_000=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_1_000=5.41e-11
.param mcrdlm4m1_cf_w_0_300_s_1_000=8.94e-12
.param mcrdlm4m1_ca_w_0_300_s_1_200=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_1_200=4.69e-11
.param mcrdlm4m1_cf_w_0_300_s_1_200=1.06e-11
.param mcrdlm4m1_ca_w_0_300_s_2_100=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_2_100=2.85e-11
.param mcrdlm4m1_cf_w_0_300_s_2_100=1.72e-11
.param mcrdlm4m1_ca_w_0_300_s_3_300=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_3_300=1.72e-11
.param mcrdlm4m1_cf_w_0_300_s_3_300=2.35e-11
.param mcrdlm4m1_ca_w_0_300_s_9_000=1.91e-05
.param mcrdlm4m1_cc_w_0_300_s_9_000=2.40e-12
.param mcrdlm4m1_cf_w_0_300_s_9_000=3.53e-11
.param mcrdlm4m1_ca_w_2_400_s_0_300=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_0_300=1.27e-10
.param mcrdlm4m1_cf_w_2_400_s_0_300=2.83e-12
.param mcrdlm4m1_ca_w_2_400_s_0_360=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_0_360=1.19e-10
.param mcrdlm4m1_cf_w_2_400_s_0_360=3.38e-12
.param mcrdlm4m1_ca_w_2_400_s_0_450=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_0_450=1.07e-10
.param mcrdlm4m1_cf_w_2_400_s_0_450=4.20e-12
.param mcrdlm4m1_ca_w_2_400_s_0_600=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_0_600=9.22e-11
.param mcrdlm4m1_cf_w_2_400_s_0_600=5.55e-12
.param mcrdlm4m1_ca_w_2_400_s_0_800=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_0_800=7.71e-11
.param mcrdlm4m1_cf_w_2_400_s_0_800=7.30e-12
.param mcrdlm4m1_ca_w_2_400_s_1_000=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_1_000=6.58e-11
.param mcrdlm4m1_cf_w_2_400_s_1_000=9.03e-12
.param mcrdlm4m1_ca_w_2_400_s_1_200=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_1_200=5.74e-11
.param mcrdlm4m1_cf_w_2_400_s_1_200=1.07e-11
.param mcrdlm4m1_ca_w_2_400_s_2_100=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_2_100=3.55e-11
.param mcrdlm4m1_cf_w_2_400_s_2_100=1.73e-11
.param mcrdlm4m1_ca_w_2_400_s_3_300=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_3_300=2.16e-11
.param mcrdlm4m1_cf_w_2_400_s_3_300=2.43e-11
.param mcrdlm4m1_ca_w_2_400_s_9_000=1.91e-05
.param mcrdlm4m1_cc_w_2_400_s_9_000=3.19e-12
.param mcrdlm4m1_cf_w_2_400_s_9_000=3.85e-11
.param mcrdlm4m2_ca_w_0_300_s_0_300=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_0_300=1.04e-10
.param mcrdlm4m2_cf_w_0_300_s_0_300=3.63e-12
.param mcrdlm4m2_ca_w_0_300_s_0_360=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_0_360=9.66e-11
.param mcrdlm4m2_cf_w_0_300_s_0_360=4.34e-12
.param mcrdlm4m2_ca_w_0_300_s_0_450=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_0_450=8.72e-11
.param mcrdlm4m2_cf_w_0_300_s_0_450=5.42e-12
.param mcrdlm4m2_ca_w_0_300_s_0_600=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_0_600=7.42e-11
.param mcrdlm4m2_cf_w_0_300_s_0_600=7.17e-12
.param mcrdlm4m2_ca_w_0_300_s_0_800=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_0_800=6.13e-11
.param mcrdlm4m2_cf_w_0_300_s_0_800=9.27e-12
.param mcrdlm4m2_ca_w_0_300_s_1_000=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_1_000=5.18e-11
.param mcrdlm4m2_cf_w_0_300_s_1_000=1.14e-11
.param mcrdlm4m2_ca_w_0_300_s_1_200=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_1_200=4.45e-11
.param mcrdlm4m2_cf_w_0_300_s_1_200=1.33e-11
.param mcrdlm4m2_ca_w_0_300_s_2_100=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_2_100=2.60e-11
.param mcrdlm4m2_cf_w_0_300_s_2_100=2.12e-11
.param mcrdlm4m2_ca_w_0_300_s_3_300=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_3_300=1.48e-11
.param mcrdlm4m2_cf_w_0_300_s_3_300=2.81e-11
.param mcrdlm4m2_ca_w_0_300_s_9_000=2.49e-05
.param mcrdlm4m2_cc_w_0_300_s_9_000=1.71e-12
.param mcrdlm4m2_cf_w_0_300_s_9_000=3.91e-11
.param mcrdlm4m2_ca_w_2_400_s_0_300=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_0_300=1.24e-10
.param mcrdlm4m2_cf_w_2_400_s_0_300=3.65e-12
.param mcrdlm4m2_ca_w_2_400_s_0_360=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_0_360=1.15e-10
.param mcrdlm4m2_cf_w_2_400_s_0_360=4.36e-12
.param mcrdlm4m2_ca_w_2_400_s_0_450=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_0_450=1.04e-10
.param mcrdlm4m2_cf_w_2_400_s_0_450=5.41e-12
.param mcrdlm4m2_ca_w_2_400_s_0_600=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_0_600=8.88e-11
.param mcrdlm4m2_cf_w_2_400_s_0_600=7.12e-12
.param mcrdlm4m2_ca_w_2_400_s_0_800=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_0_800=7.37e-11
.param mcrdlm4m2_cf_w_2_400_s_0_800=9.33e-12
.param mcrdlm4m2_ca_w_2_400_s_1_000=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_1_000=6.26e-11
.param mcrdlm4m2_cf_w_2_400_s_1_000=1.15e-11
.param mcrdlm4m2_ca_w_2_400_s_1_200=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_1_200=5.40e-11
.param mcrdlm4m2_cf_w_2_400_s_1_200=1.35e-11
.param mcrdlm4m2_ca_w_2_400_s_2_100=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_2_100=3.24e-11
.param mcrdlm4m2_cf_w_2_400_s_2_100=2.14e-11
.param mcrdlm4m2_ca_w_2_400_s_3_300=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_3_300=1.89e-11
.param mcrdlm4m2_cf_w_2_400_s_3_300=2.91e-11
.param mcrdlm4m2_ca_w_2_400_s_9_000=2.49e-05
.param mcrdlm4m2_cc_w_2_400_s_9_000=2.37e-12
.param mcrdlm4m2_cf_w_2_400_s_9_000=4.26e-11
.param mcrdlm4m3_ca_w_0_300_s_0_300=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_0_300=9.29e-11
.param mcrdlm4m3_cf_w_0_300_s_0_300=1.24e-11
.param mcrdlm4m3_ca_w_0_300_s_0_360=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_0_360=8.49e-11
.param mcrdlm4m3_cf_w_0_300_s_0_360=1.46e-11
.param mcrdlm4m3_ca_w_0_300_s_0_450=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_0_450=7.50e-11
.param mcrdlm4m3_cf_w_0_300_s_0_450=1.77e-11
.param mcrdlm4m3_ca_w_0_300_s_0_600=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_0_600=6.16e-11
.param mcrdlm4m3_cf_w_0_300_s_0_600=2.23e-11
.param mcrdlm4m3_ca_w_0_300_s_0_800=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_0_800=4.89e-11
.param mcrdlm4m3_cf_w_0_300_s_0_800=2.74e-11
.param mcrdlm4m3_ca_w_0_300_s_1_000=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_1_000=3.94e-11
.param mcrdlm4m3_cf_w_0_300_s_1_000=3.19e-11
.param mcrdlm4m3_ca_w_0_300_s_1_200=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_1_200=3.23e-11
.param mcrdlm4m3_cf_w_0_300_s_1_200=3.56e-11
.param mcrdlm4m3_ca_w_0_300_s_2_100=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_2_100=1.56e-11
.param mcrdlm4m3_cf_w_0_300_s_2_100=4.70e-11
.param mcrdlm4m3_ca_w_0_300_s_3_300=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_3_300=7.52e-12
.param mcrdlm4m3_cf_w_0_300_s_3_300=5.39e-11
.param mcrdlm4m3_ca_w_0_300_s_9_000=9.25e-05
.param mcrdlm4m3_cc_w_0_300_s_9_000=5.95e-13
.param mcrdlm4m3_cf_w_0_300_s_9_000=6.04e-11
.param mcrdlm4m3_ca_w_2_400_s_0_300=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_0_300=1.09e-10
.param mcrdlm4m3_cf_w_2_400_s_0_300=1.24e-11
.param mcrdlm4m3_ca_w_2_400_s_0_360=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_0_360=9.95e-11
.param mcrdlm4m3_cf_w_2_400_s_0_360=1.46e-11
.param mcrdlm4m3_ca_w_2_400_s_0_450=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_0_450=8.85e-11
.param mcrdlm4m3_cf_w_2_400_s_0_450=1.77e-11
.param mcrdlm4m3_ca_w_2_400_s_0_600=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_0_600=7.37e-11
.param mcrdlm4m3_cf_w_2_400_s_0_600=2.23e-11
.param mcrdlm4m3_ca_w_2_400_s_0_800=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_0_800=5.92e-11
.param mcrdlm4m3_cf_w_2_400_s_0_800=2.75e-11
.param mcrdlm4m3_ca_w_2_400_s_1_000=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_1_000=4.84e-11
.param mcrdlm4m3_cf_w_2_400_s_1_000=3.20e-11
.param mcrdlm4m3_ca_w_2_400_s_1_200=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_1_200=4.06e-11
.param mcrdlm4m3_cf_w_2_400_s_1_200=3.58e-11
.param mcrdlm4m3_ca_w_2_400_s_2_100=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_2_100=2.16e-11
.param mcrdlm4m3_cf_w_2_400_s_2_100=4.75e-11
.param mcrdlm4m3_ca_w_2_400_s_3_300=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_3_300=1.11e-11
.param mcrdlm4m3_cf_w_2_400_s_3_300=5.59e-11
.param mcrdlm4m3_ca_w_2_400_s_9_000=9.25e-05
.param mcrdlm4m3_cc_w_2_400_s_9_000=9.05e-13
.param mcrdlm4m3_cf_w_2_400_s_9_000=6.53e-11
.param mcrdlm5f_ca_w_1_600_s_1_600=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_1_600=6.69e-11
.param mcrdlm5f_cf_w_1_600_s_1_600=9.13e-12
.param mcrdlm5f_ca_w_1_600_s_1_700=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_1_700=6.30e-11
.param mcrdlm5f_cf_w_1_600_s_1_700=9.67e-12
.param mcrdlm5f_ca_w_1_600_s_1_900=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_1_900=5.65e-11
.param mcrdlm5f_cf_w_1_600_s_1_900=1.07e-11
.param mcrdlm5f_ca_w_1_600_s_2_000=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_2_000=5.37e-11
.param mcrdlm5f_cf_w_1_600_s_2_000=1.12e-11
.param mcrdlm5f_ca_w_1_600_s_2_400=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_2_400=4.48e-11
.param mcrdlm5f_cf_w_1_600_s_2_400=1.33e-11
.param mcrdlm5f_ca_w_1_600_s_2_800=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_2_800=3.82e-11
.param mcrdlm5f_cf_w_1_600_s_2_800=1.52e-11
.param mcrdlm5f_ca_w_1_600_s_3_200=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_3_200=3.30e-11
.param mcrdlm5f_cf_w_1_600_s_3_200=1.70e-11
.param mcrdlm5f_ca_w_1_600_s_4_800=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_4_800=1.99e-11
.param mcrdlm5f_cf_w_1_600_s_4_800=2.33e-11
.param mcrdlm5f_ca_w_1_600_s_10_000=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_10_000=4.80e-12
.param mcrdlm5f_cf_w_1_600_s_10_000=3.43e-11
.param mcrdlm5f_ca_w_1_600_s_12_000=1.20e-05
.param mcrdlm5f_cc_w_1_600_s_12_000=2.83e-12
.param mcrdlm5f_cf_w_1_600_s_12_000=3.61e-11
.param mcrdlm5f_ca_w_4_000_s_1_600=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_1_600=6.99e-11
.param mcrdlm5f_cf_w_4_000_s_1_600=9.13e-12
.param mcrdlm5f_ca_w_4_000_s_1_700=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_1_700=6.59e-11
.param mcrdlm5f_cf_w_4_000_s_1_700=9.67e-12
.param mcrdlm5f_ca_w_4_000_s_1_900=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_1_900=5.91e-11
.param mcrdlm5f_cf_w_4_000_s_1_900=1.07e-11
.param mcrdlm5f_ca_w_4_000_s_2_000=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_2_000=5.62e-11
.param mcrdlm5f_cf_w_4_000_s_2_000=1.13e-11
.param mcrdlm5f_ca_w_4_000_s_2_400=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_2_400=4.69e-11
.param mcrdlm5f_cf_w_4_000_s_2_400=1.33e-11
.param mcrdlm5f_ca_w_4_000_s_2_800=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_2_800=4.00e-11
.param mcrdlm5f_cf_w_4_000_s_2_800=1.52e-11
.param mcrdlm5f_ca_w_4_000_s_3_200=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_3_200=3.47e-11
.param mcrdlm5f_cf_w_4_000_s_3_200=1.71e-11
.param mcrdlm5f_ca_w_4_000_s_4_800=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_4_800=2.09e-11
.param mcrdlm5f_cf_w_4_000_s_4_800=2.35e-11
.param mcrdlm5f_ca_w_4_000_s_10_000=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_10_000=5.08e-12
.param mcrdlm5f_cf_w_4_000_s_10_000=3.49e-11
.param mcrdlm5f_ca_w_4_000_s_12_000=1.20e-05
.param mcrdlm5f_cc_w_4_000_s_12_000=3.03e-12
.param mcrdlm5f_cf_w_4_000_s_12_000=3.68e-11
.param mcrdlm5d_ca_w_1_600_s_1_600=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_1_600=6.64e-11
.param mcrdlm5d_cf_w_1_600_s_1_600=9.43e-12
.param mcrdlm5d_ca_w_1_600_s_1_700=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_1_700=6.25e-11
.param mcrdlm5d_cf_w_1_600_s_1_700=9.98e-12
.param mcrdlm5d_ca_w_1_600_s_1_900=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_1_900=5.60e-11
.param mcrdlm5d_cf_w_1_600_s_1_900=1.11e-11
.param mcrdlm5d_ca_w_1_600_s_2_000=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_2_000=5.32e-11
.param mcrdlm5d_cf_w_1_600_s_2_000=1.16e-11
.param mcrdlm5d_ca_w_1_600_s_2_400=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_2_400=4.42e-11
.param mcrdlm5d_cf_w_1_600_s_2_400=1.37e-11
.param mcrdlm5d_ca_w_1_600_s_2_800=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_2_800=3.77e-11
.param mcrdlm5d_cf_w_1_600_s_2_800=1.57e-11
.param mcrdlm5d_ca_w_1_600_s_3_200=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_3_200=3.25e-11
.param mcrdlm5d_cf_w_1_600_s_3_200=1.76e-11
.param mcrdlm5d_ca_w_1_600_s_4_800=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_4_800=1.94e-11
.param mcrdlm5d_cf_w_1_600_s_4_800=2.40e-11
.param mcrdlm5d_ca_w_1_600_s_10_000=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_10_000=4.51e-12
.param mcrdlm5d_cf_w_1_600_s_10_000=3.49e-11
.param mcrdlm5d_ca_w_1_600_s_12_000=1.24e-05
.param mcrdlm5d_cc_w_1_600_s_12_000=2.62e-12
.param mcrdlm5d_cf_w_1_600_s_12_000=3.66e-11
.param mcrdlm5d_ca_w_4_000_s_1_600=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_1_600=6.93e-11
.param mcrdlm5d_cf_w_4_000_s_1_600=9.42e-12
.param mcrdlm5d_ca_w_4_000_s_1_700=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_1_700=6.54e-11
.param mcrdlm5d_cf_w_4_000_s_1_700=9.98e-12
.param mcrdlm5d_ca_w_4_000_s_1_900=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_1_900=5.86e-11
.param mcrdlm5d_cf_w_4_000_s_1_900=1.11e-11
.param mcrdlm5d_ca_w_4_000_s_2_000=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_2_000=5.57e-11
.param mcrdlm5d_cf_w_4_000_s_2_000=1.16e-11
.param mcrdlm5d_ca_w_4_000_s_2_400=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_2_400=4.63e-11
.param mcrdlm5d_cf_w_4_000_s_2_400=1.37e-11
.param mcrdlm5d_ca_w_4_000_s_2_800=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_2_800=3.94e-11
.param mcrdlm5d_cf_w_4_000_s_2_800=1.57e-11
.param mcrdlm5d_ca_w_4_000_s_3_200=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_3_200=3.40e-11
.param mcrdlm5d_cf_w_4_000_s_3_200=1.76e-11
.param mcrdlm5d_ca_w_4_000_s_4_800=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_4_800=2.03e-11
.param mcrdlm5d_cf_w_4_000_s_4_800=2.41e-11
.param mcrdlm5d_ca_w_4_000_s_10_000=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_10_000=4.75e-12
.param mcrdlm5d_cf_w_4_000_s_10_000=3.55e-11
.param mcrdlm5d_ca_w_4_000_s_12_000=1.24e-05
.param mcrdlm5d_cc_w_4_000_s_12_000=2.79e-12
.param mcrdlm5d_cf_w_4_000_s_12_000=3.73e-11
.param mcrdlm5p1_ca_w_1_600_s_1_600=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_1_600=6.60e-11
.param mcrdlm5p1_cf_w_1_600_s_1_600=9.71e-12
.param mcrdlm5p1_ca_w_1_600_s_1_700=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_1_700=6.21e-11
.param mcrdlm5p1_cf_w_1_600_s_1_700=1.03e-11
.param mcrdlm5p1_ca_w_1_600_s_1_900=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_1_900=5.57e-11
.param mcrdlm5p1_cf_w_1_600_s_1_900=1.14e-11
.param mcrdlm5p1_ca_w_1_600_s_2_000=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_2_000=5.29e-11
.param mcrdlm5p1_cf_w_1_600_s_2_000=1.19e-11
.param mcrdlm5p1_ca_w_1_600_s_2_400=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_2_400=4.38e-11
.param mcrdlm5p1_cf_w_1_600_s_2_400=1.41e-11
.param mcrdlm5p1_ca_w_1_600_s_2_800=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_2_800=3.73e-11
.param mcrdlm5p1_cf_w_1_600_s_2_800=1.61e-11
.param mcrdlm5p1_ca_w_1_600_s_3_200=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_3_200=3.21e-11
.param mcrdlm5p1_cf_w_1_600_s_3_200=1.81e-11
.param mcrdlm5p1_ca_w_1_600_s_4_800=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_4_800=1.90e-11
.param mcrdlm5p1_cf_w_1_600_s_4_800=2.46e-11
.param mcrdlm5p1_ca_w_1_600_s_10_000=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_10_000=4.25e-12
.param mcrdlm5p1_cf_w_1_600_s_10_000=3.55e-11
.param mcrdlm5p1_ca_w_1_600_s_12_000=1.27e-05
.param mcrdlm5p1_cc_w_1_600_s_12_000=2.44e-12
.param mcrdlm5p1_cf_w_1_600_s_12_000=3.72e-11
.param mcrdlm5p1_ca_w_4_000_s_1_600=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_1_600=6.88e-11
.param mcrdlm5p1_cf_w_4_000_s_1_600=9.71e-12
.param mcrdlm5p1_ca_w_4_000_s_1_700=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_1_700=6.47e-11
.param mcrdlm5p1_cf_w_4_000_s_1_700=1.03e-11
.param mcrdlm5p1_ca_w_4_000_s_1_900=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_1_900=5.80e-11
.param mcrdlm5p1_cf_w_4_000_s_1_900=1.14e-11
.param mcrdlm5p1_ca_w_4_000_s_2_000=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_2_000=5.51e-11
.param mcrdlm5p1_cf_w_4_000_s_2_000=1.20e-11
.param mcrdlm5p1_ca_w_4_000_s_2_400=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_2_400=4.59e-11
.param mcrdlm5p1_cf_w_4_000_s_2_400=1.41e-11
.param mcrdlm5p1_ca_w_4_000_s_2_800=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_2_800=3.89e-11
.param mcrdlm5p1_cf_w_4_000_s_2_800=1.62e-11
.param mcrdlm5p1_ca_w_4_000_s_3_200=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_3_200=3.35e-11
.param mcrdlm5p1_cf_w_4_000_s_3_200=1.81e-11
.param mcrdlm5p1_ca_w_4_000_s_4_800=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_4_800=1.98e-11
.param mcrdlm5p1_cf_w_4_000_s_4_800=2.47e-11
.param mcrdlm5p1_ca_w_4_000_s_10_000=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_10_000=4.47e-12
.param mcrdlm5p1_cf_w_4_000_s_10_000=3.61e-11
.param mcrdlm5p1_ca_w_4_000_s_12_000=1.27e-05
.param mcrdlm5p1_cc_w_4_000_s_12_000=2.57e-12
.param mcrdlm5p1_cf_w_4_000_s_12_000=3.79e-11
.param mcrdlm5l1_ca_w_1_600_s_1_600=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_1_600=6.52e-11
.param mcrdlm5l1_cf_w_1_600_s_1_600=1.03e-11
.param mcrdlm5l1_ca_w_1_600_s_1_700=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_1_700=6.13e-11
.param mcrdlm5l1_cf_w_1_600_s_1_700=1.09e-11
.param mcrdlm5l1_ca_w_1_600_s_1_900=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_1_900=5.49e-11
.param mcrdlm5l1_cf_w_1_600_s_1_900=1.20e-11
.param mcrdlm5l1_ca_w_1_600_s_2_000=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_2_000=5.21e-11
.param mcrdlm5l1_cf_w_1_600_s_2_000=1.26e-11
.param mcrdlm5l1_ca_w_1_600_s_2_400=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_2_400=4.30e-11
.param mcrdlm5l1_cf_w_1_600_s_2_400=1.49e-11
.param mcrdlm5l1_ca_w_1_600_s_2_800=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_2_800=3.64e-11
.param mcrdlm5l1_cf_w_1_600_s_2_800=1.70e-11
.param mcrdlm5l1_ca_w_1_600_s_3_200=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_3_200=3.12e-11
.param mcrdlm5l1_cf_w_1_600_s_3_200=1.90e-11
.param mcrdlm5l1_ca_w_1_600_s_4_800=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_4_800=1.81e-11
.param mcrdlm5l1_cf_w_1_600_s_4_800=2.58e-11
.param mcrdlm5l1_ca_w_1_600_s_10_000=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_10_000=3.79e-12
.param mcrdlm5l1_cf_w_1_600_s_10_000=3.66e-11
.param mcrdlm5l1_ca_w_1_600_s_12_000=1.35e-05
.param mcrdlm5l1_cc_w_1_600_s_12_000=2.14e-12
.param mcrdlm5l1_cf_w_1_600_s_12_000=3.82e-11
.param mcrdlm5l1_ca_w_4_000_s_1_600=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_1_600=6.77e-11
.param mcrdlm5l1_cf_w_4_000_s_1_600=1.03e-11
.param mcrdlm5l1_ca_w_4_000_s_1_700=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_1_700=6.37e-11
.param mcrdlm5l1_cf_w_4_000_s_1_700=1.09e-11
.param mcrdlm5l1_ca_w_4_000_s_1_900=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_1_900=5.70e-11
.param mcrdlm5l1_cf_w_4_000_s_1_900=1.21e-11
.param mcrdlm5l1_ca_w_4_000_s_2_000=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_2_000=5.41e-11
.param mcrdlm5l1_cf_w_4_000_s_2_000=1.26e-11
.param mcrdlm5l1_ca_w_4_000_s_2_400=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_2_400=4.48e-11
.param mcrdlm5l1_cf_w_4_000_s_2_400=1.49e-11
.param mcrdlm5l1_ca_w_4_000_s_2_800=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_2_800=3.78e-11
.param mcrdlm5l1_cf_w_4_000_s_2_800=1.70e-11
.param mcrdlm5l1_ca_w_4_000_s_3_200=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_3_200=3.25e-11
.param mcrdlm5l1_cf_w_4_000_s_3_200=1.91e-11
.param mcrdlm5l1_ca_w_4_000_s_4_800=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_4_800=1.89e-11
.param mcrdlm5l1_cf_w_4_000_s_4_800=2.59e-11
.param mcrdlm5l1_ca_w_4_000_s_10_000=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_10_000=4.01e-12
.param mcrdlm5l1_cf_w_4_000_s_10_000=3.72e-11
.param mcrdlm5l1_ca_w_4_000_s_12_000=1.35e-05
.param mcrdlm5l1_cc_w_4_000_s_12_000=2.28e-12
.param mcrdlm5l1_cf_w_4_000_s_12_000=3.89e-11
.param mcrdlm5m1_ca_w_1_600_s_1_600=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_1_600=6.39e-11
.param mcrdlm5m1_cf_w_1_600_s_1_600=1.13e-11
.param mcrdlm5m1_ca_w_1_600_s_1_700=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_1_700=5.99e-11
.param mcrdlm5m1_cf_w_1_600_s_1_700=1.20e-11
.param mcrdlm5m1_ca_w_1_600_s_1_900=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_1_900=5.35e-11
.param mcrdlm5m1_cf_w_1_600_s_1_900=1.33e-11
.param mcrdlm5m1_ca_w_1_600_s_2_000=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_2_000=5.06e-11
.param mcrdlm5m1_cf_w_1_600_s_2_000=1.39e-11
.param mcrdlm5m1_ca_w_1_600_s_2_400=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_2_400=4.15e-11
.param mcrdlm5m1_cf_w_1_600_s_2_400=1.63e-11
.param mcrdlm5m1_ca_w_1_600_s_2_800=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_2_800=3.49e-11
.param mcrdlm5m1_cf_w_1_600_s_2_800=1.86e-11
.param mcrdlm5m1_ca_w_1_600_s_3_200=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_3_200=2.97e-11
.param mcrdlm5m1_cf_w_1_600_s_3_200=2.08e-11
.param mcrdlm5m1_ca_w_1_600_s_4_800=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_4_800=1.67e-11
.param mcrdlm5m1_cf_w_1_600_s_4_800=2.79e-11
.param mcrdlm5m1_ca_w_1_600_s_10_000=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_10_000=3.12e-12
.param mcrdlm5m1_cf_w_1_600_s_10_000=3.85e-11
.param mcrdlm5m1_ca_w_1_600_s_12_000=1.50e-05
.param mcrdlm5m1_cc_w_1_600_s_12_000=1.66e-12
.param mcrdlm5m1_cf_w_1_600_s_12_000=4.00e-11
.param mcrdlm5m1_ca_w_4_000_s_1_600=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_1_600=6.60e-11
.param mcrdlm5m1_cf_w_4_000_s_1_600=1.13e-11
.param mcrdlm5m1_ca_w_4_000_s_1_700=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_1_700=6.21e-11
.param mcrdlm5m1_cf_w_4_000_s_1_700=1.20e-11
.param mcrdlm5m1_ca_w_4_000_s_1_900=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_1_900=5.53e-11
.param mcrdlm5m1_cf_w_4_000_s_1_900=1.33e-11
.param mcrdlm5m1_ca_w_4_000_s_2_000=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_2_000=5.24e-11
.param mcrdlm5m1_cf_w_4_000_s_2_000=1.39e-11
.param mcrdlm5m1_ca_w_4_000_s_2_400=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_2_400=4.32e-11
.param mcrdlm5m1_cf_w_4_000_s_2_400=1.64e-11
.param mcrdlm5m1_ca_w_4_000_s_2_800=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_2_800=3.61e-11
.param mcrdlm5m1_cf_w_4_000_s_2_800=1.87e-11
.param mcrdlm5m1_ca_w_4_000_s_3_200=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_3_200=3.07e-11
.param mcrdlm5m1_cf_w_4_000_s_3_200=2.09e-11
.param mcrdlm5m1_ca_w_4_000_s_4_800=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_4_800=1.74e-11
.param mcrdlm5m1_cf_w_4_000_s_4_800=2.81e-11
.param mcrdlm5m1_ca_w_4_000_s_10_000=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_10_000=3.30e-12
.param mcrdlm5m1_cf_w_4_000_s_10_000=3.91e-11
.param mcrdlm5m1_ca_w_4_000_s_12_000=1.50e-05
.param mcrdlm5m1_cc_w_4_000_s_12_000=1.76e-12
.param mcrdlm5m1_cf_w_4_000_s_12_000=4.06e-11
.param mcrdlm5m2_ca_w_1_600_s_1_600=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_1_600=6.22e-11
.param mcrdlm5m2_cf_w_1_600_s_1_600=1.27e-11
.param mcrdlm5m2_ca_w_1_600_s_1_700=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_1_700=5.83e-11
.param mcrdlm5m2_cf_w_1_600_s_1_700=1.35e-11
.param mcrdlm5m2_ca_w_1_600_s_1_900=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_1_900=5.17e-11
.param mcrdlm5m2_cf_w_1_600_s_1_900=1.49e-11
.param mcrdlm5m2_ca_w_1_600_s_2_000=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_2_000=4.88e-11
.param mcrdlm5m2_cf_w_1_600_s_2_000=1.56e-11
.param mcrdlm5m2_ca_w_1_600_s_2_400=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_2_400=3.98e-11
.param mcrdlm5m2_cf_w_1_600_s_2_400=1.83e-11
.param mcrdlm5m2_ca_w_1_600_s_2_800=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_2_800=3.31e-11
.param mcrdlm5m2_cf_w_1_600_s_2_800=2.08e-11
.param mcrdlm5m2_ca_w_1_600_s_3_200=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_3_200=2.79e-11
.param mcrdlm5m2_cf_w_1_600_s_3_200=2.31e-11
.param mcrdlm5m2_ca_w_1_600_s_4_800=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_4_800=1.51e-11
.param mcrdlm5m2_cf_w_1_600_s_4_800=3.06e-11
.param mcrdlm5m2_ca_w_1_600_s_10_000=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_10_000=2.48e-12
.param mcrdlm5m2_cf_w_1_600_s_10_000=4.09e-11
.param mcrdlm5m2_ca_w_1_600_s_12_000=1.70e-05
.param mcrdlm5m2_cc_w_1_600_s_12_000=1.27e-12
.param mcrdlm5m2_cf_w_1_600_s_12_000=4.21e-11
.param mcrdlm5m2_ca_w_4_000_s_1_600=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_1_600=6.41e-11
.param mcrdlm5m2_cf_w_4_000_s_1_600=1.27e-11
.param mcrdlm5m2_ca_w_4_000_s_1_700=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_1_700=6.01e-11
.param mcrdlm5m2_cf_w_4_000_s_1_700=1.35e-11
.param mcrdlm5m2_ca_w_4_000_s_1_900=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_1_900=5.33e-11
.param mcrdlm5m2_cf_w_4_000_s_1_900=1.49e-11
.param mcrdlm5m2_ca_w_4_000_s_2_000=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_2_000=5.03e-11
.param mcrdlm5m2_cf_w_4_000_s_2_000=1.56e-11
.param mcrdlm5m2_ca_w_4_000_s_2_400=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_2_400=4.11e-11
.param mcrdlm5m2_cf_w_4_000_s_2_400=1.83e-11
.param mcrdlm5m2_ca_w_4_000_s_2_800=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_2_800=3.42e-11
.param mcrdlm5m2_cf_w_4_000_s_2_800=2.08e-11
.param mcrdlm5m2_ca_w_4_000_s_3_200=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_3_200=2.89e-11
.param mcrdlm5m2_cf_w_4_000_s_3_200=2.32e-11
.param mcrdlm5m2_ca_w_4_000_s_4_800=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_4_800=1.57e-11
.param mcrdlm5m2_cf_w_4_000_s_4_800=3.08e-11
.param mcrdlm5m2_ca_w_4_000_s_10_000=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_10_000=2.60e-12
.param mcrdlm5m2_cf_w_4_000_s_10_000=4.14e-11
.param mcrdlm5m2_ca_w_4_000_s_12_000=1.70e-05
.param mcrdlm5m2_cc_w_4_000_s_12_000=1.32e-12
.param mcrdlm5m2_cf_w_4_000_s_12_000=4.27e-11
.param mcrdlm5m3_ca_w_1_600_s_1_600=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_1_600=5.67e-11
.param mcrdlm5m3_cf_w_1_600_s_1_600=1.83e-11
.param mcrdlm5m3_ca_w_1_600_s_1_700=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_1_700=5.28e-11
.param mcrdlm5m3_cf_w_1_600_s_1_700=1.93e-11
.param mcrdlm5m3_ca_w_1_600_s_1_900=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_1_900=4.62e-11
.param mcrdlm5m3_cf_w_1_600_s_1_900=2.12e-11
.param mcrdlm5m3_ca_w_1_600_s_2_000=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_2_000=4.34e-11
.param mcrdlm5m3_cf_w_1_600_s_2_000=2.22e-11
.param mcrdlm5m3_ca_w_1_600_s_2_400=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_2_400=3.44e-11
.param mcrdlm5m3_cf_w_1_600_s_2_400=2.57e-11
.param mcrdlm5m3_ca_w_1_600_s_2_800=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_2_800=2.79e-11
.param mcrdlm5m3_cf_w_1_600_s_2_800=2.88e-11
.param mcrdlm5m3_ca_w_1_600_s_3_200=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_3_200=2.29e-11
.param mcrdlm5m3_cf_w_1_600_s_3_200=3.16e-11
.param mcrdlm5m3_ca_w_1_600_s_4_800=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_4_800=1.10e-11
.param mcrdlm5m3_cf_w_1_600_s_4_800=3.98e-11
.param mcrdlm5m3_ca_w_1_600_s_10_000=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_10_000=1.26e-12
.param mcrdlm5m3_cf_w_1_600_s_10_000=4.85e-11
.param mcrdlm5m3_ca_w_1_600_s_12_000=2.53e-05
.param mcrdlm5m3_cc_w_1_600_s_12_000=5.70e-13
.param mcrdlm5m3_cf_w_1_600_s_12_000=4.92e-11
.param mcrdlm5m3_ca_w_4_000_s_1_600=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_1_600=5.82e-11
.param mcrdlm5m3_cf_w_4_000_s_1_600=1.83e-11
.param mcrdlm5m3_ca_w_4_000_s_1_700=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_1_700=5.42e-11
.param mcrdlm5m3_cf_w_4_000_s_1_700=1.93e-11
.param mcrdlm5m3_ca_w_4_000_s_1_900=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_1_900=4.75e-11
.param mcrdlm5m3_cf_w_4_000_s_1_900=2.12e-11
.param mcrdlm5m3_ca_w_4_000_s_2_000=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_2_000=4.46e-11
.param mcrdlm5m3_cf_w_4_000_s_2_000=2.22e-11
.param mcrdlm5m3_ca_w_4_000_s_2_400=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_2_400=3.53e-11
.param mcrdlm5m3_cf_w_4_000_s_2_400=2.57e-11
.param mcrdlm5m3_ca_w_4_000_s_2_800=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_2_800=2.87e-11
.param mcrdlm5m3_cf_w_4_000_s_2_800=2.89e-11
.param mcrdlm5m3_ca_w_4_000_s_3_200=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_3_200=2.36e-11
.param mcrdlm5m3_cf_w_4_000_s_3_200=3.17e-11
.param mcrdlm5m3_ca_w_4_000_s_4_800=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_4_800=1.14e-11
.param mcrdlm5m3_cf_w_4_000_s_4_800=4.00e-11
.param mcrdlm5m3_ca_w_4_000_s_10_000=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_10_000=1.33e-12
.param mcrdlm5m3_cf_w_4_000_s_10_000=4.90e-11
.param mcrdlm5m3_ca_w_4_000_s_12_000=2.53e-05
.param mcrdlm5m3_cc_w_4_000_s_12_000=6.30e-13
.param mcrdlm5m3_cf_w_4_000_s_12_000=4.97e-11
.param mcrdlm5m4_ca_w_1_600_s_1_600=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_1_600=4.40e-11
.param mcrdlm5m4_cf_w_1_600_s_1_600=4.21e-11
.param mcrdlm5m4_ca_w_1_600_s_1_700=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_1_700=4.03e-11
.param mcrdlm5m4_cf_w_1_600_s_1_700=4.38e-11
.param mcrdlm5m4_ca_w_1_600_s_1_900=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_1_900=3.40e-11
.param mcrdlm5m4_cf_w_1_600_s_1_900=4.70e-11
.param mcrdlm5m4_ca_w_1_600_s_2_000=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_2_000=3.15e-11
.param mcrdlm5m4_cf_w_1_600_s_2_000=4.84e-11
.param mcrdlm5m4_ca_w_1_600_s_2_400=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_2_400=2.33e-11
.param mcrdlm5m4_cf_w_1_600_s_2_400=5.34e-11
.param mcrdlm5m4_ca_w_1_600_s_2_800=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_2_800=1.77e-11
.param mcrdlm5m4_cf_w_1_600_s_2_800=5.73e-11
.param mcrdlm5m4_ca_w_1_600_s_3_200=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_3_200=1.37e-11
.param mcrdlm5m4_cf_w_1_600_s_3_200=6.03e-11
.param mcrdlm5m4_ca_w_1_600_s_4_800=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_4_800=5.39e-12
.param mcrdlm5m4_cf_w_1_600_s_4_800=6.74e-11
.param mcrdlm5m4_ca_w_1_600_s_10_000=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_10_000=4.30e-13
.param mcrdlm5m4_cf_w_1_600_s_10_000=7.23e-11
.param mcrdlm5m4_ca_w_1_600_s_12_000=7.39e-05
.param mcrdlm5m4_cc_w_1_600_s_12_000=1.80e-13
.param mcrdlm5m4_cf_w_1_600_s_12_000=7.25e-11
.param mcrdlm5m4_ca_w_4_000_s_1_600=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_1_600=4.55e-11
.param mcrdlm5m4_cf_w_4_000_s_1_600=4.22e-11
.param mcrdlm5m4_ca_w_4_000_s_1_700=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_1_700=4.16e-11
.param mcrdlm5m4_cf_w_4_000_s_1_700=4.39e-11
.param mcrdlm5m4_ca_w_4_000_s_1_900=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_1_900=3.53e-11
.param mcrdlm5m4_cf_w_4_000_s_1_900=4.70e-11
.param mcrdlm5m4_ca_w_4_000_s_2_000=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_2_000=3.25e-11
.param mcrdlm5m4_cf_w_4_000_s_2_000=4.83e-11
.param mcrdlm5m4_ca_w_4_000_s_2_400=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_2_400=2.43e-11
.param mcrdlm5m4_cf_w_4_000_s_2_400=5.33e-11
.param mcrdlm5m4_ca_w_4_000_s_2_800=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_2_800=1.86e-11
.param mcrdlm5m4_cf_w_4_000_s_2_800=5.73e-11
.param mcrdlm5m4_ca_w_4_000_s_3_200=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_3_200=1.44e-11
.param mcrdlm5m4_cf_w_4_000_s_3_200=6.05e-11
.param mcrdlm5m4_ca_w_4_000_s_4_800=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_4_800=5.85e-12
.param mcrdlm5m4_cf_w_4_000_s_4_800=6.77e-11
.param mcrdlm5m4_ca_w_4_000_s_10_000=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_10_000=4.45e-13
.param mcrdlm5m4_cf_w_4_000_s_10_000=7.29e-11
.param mcrdlm5m4_ca_w_4_000_s_12_000=7.39e-05
.param mcrdlm5m4_cc_w_4_000_s_12_000=1.80e-13
.param mcrdlm5m4_cf_w_4_000_s_12_000=7.32e-11
.param cp1f=1.06e-04
.param cp1fsw=8.64e-11
.param cl1f=3.69e-05
.param cl1fsw=8.30e-11
.param cl1d=5.53e-05
.param cl1dsw=8.23e-11
.param cl1p1=9.41e-05
.param cl1p1sw=8.13e-11
.param cm1f=2.58e-05
.param cm1fsw=1.07e-10
.param cm1d=3.36e-05
.param cm1dsw=1.06e-10
.param cm1p1=4.48e-05
.param cm1p1sw=1.06e-10
.param cm1l1=1.14e-04
.param cm1l1sw=1.03e-10
.param cm2f=1.75e-05
.param cm2fsw=1.08e-10
.param cm2d=2.08e-05
.param cm2dsw=1.07e-10
.param cm2p1=2.47e-05
.param cm2p1sw=1.07e-10
.param cm2l1=3.70e-05
.param cm2l1sw=1.06e-10
.param cm2m1=1.28e-04
.param cm2m1sw=1.03e-10
.param cm3f=1.26e-05
.param cm3fsw=1.08e-10
.param cm3d=1.42e-05
.param cm3dsw=1.09e-10
.param cm3p1=1.58e-05
.param cm3p1sw=1.08e-10
.param cm3l1=2.02e-05
.param cm3l1sw=1.08e-10
.param cm3m1=3.29e-05
.param cm3m1sw=1.07e-10
.param cm3m2=8.22e-05
.param cm3m2sw=1.05e-10
.param cm4f=8.67e-06
.param cm4fsw=1.09e-10
.param cm4d=9.41e-06
.param cm4dsw=1.09e-10
.param cm4p1=1.01e-05
.param cm4p1sw=1.09e-10
.param cm4l1=1.17e-05
.param cm4l1sw=1.09e-10
.param cm4m1=1.51e-05
.param cm4m1sw=1.08e-10
.param cm4m2=2.09e-05
.param cm4m2sw=1.08e-10
.param cm4m3=8.85e-05
.param cm4m3sw=1.05e-10
.param cm5f=6.48e-06
.param cm5fsw=7.85e-11
.param cm5d=6.88e-06
.param cm5dsw=7.84e-11
.param cm5p1=7.26e-06
.param cm5p1sw=7.82e-11
.param cm5l1=8.04e-06
.param cm5l1sw=7.80e-11
.param cm5m1=9.50e-06
.param cm5m1sw=7.77e-11
.param cm5m2=1.15e-05
.param cm5m2sw=7.74e-11
.param cm5m3=1.99e-05
.param cm5m3sw=7.76e-11
.param cm5m4=6.84e-05
.param cm5m4sw=8.87e-11
.param crdlf=2.57e-06
.param crdlfsw=5.75e-11
.param crdld=2.63e-06
.param crdldsw=5.75e-11
.param crdlp1=2.68e-06
.param crdlp1sw=5.74e-11
.param crdll1=2.78e-06
.param crdll1sw=5.73e-11
.param crdlm1=2.93e-06
.param crdlm1sw=5.71e-11
.param crdlm2=3.10e-06
.param crdlm2sw=5.70e-11
.param crdlm3=3.50e-06
.param crdlm3sw=5.68e-11
.param crdlm4=4.00e-06
.param crdlm4sw=5.66e-11
.param crdlm5=5.44e-06
.param crdlm5sw=5.68e-11
.param cl1p1f=2.00e-04
.param cl1p1fsw=8.32e-11
.param cm1p1f=1.51e-04
.param cm1p1fsw=8.45e-11
.param cm2p1f=1.31e-04
.param cm2p1fsw=8.53e-11
.param cm3p1f=1.22e-04
.param cm3p1fsw=8.58e-11
.param cm4p1f=1.16e-04
.param cm4p1fsw=8.61e-11
.param cm5p1f=1.13e-04
.param cm5p1fsw=8.61e-11
.param crdlp1f=1.09e-04
.param crdlp1fsw=8.63e-11
.param cm1l1f=1.51e-04
.param cm1l1fsw=7.90e-11
.param cm1l1d=1.69e-04
.param cm1l1dsw=7.81e-11
.param cm1l1p1=2.08e-04
.param cm1l1p1sw=7.71e-11
.param cm2l1f=7.40e-05
.param cm2l1fsw=8.14e-11
.param cm2l1d=9.23e-05
.param cm2l1dsw=8.04e-11
.param cm2l1p1=1.31e-04
.param cm2l1p1sw=7.94e-11
.param cm3l1f=5.71e-05
.param cm3l1fsw=8.21e-11
.param cm3l1d=7.54e-05
.param cm3l1dsw=8.13e-11
.param cm3l1p1=1.14e-04
.param cm3l1p1sw=8.04e-11
.param cm4l1f=4.86e-05
.param cm4l1fsw=8.26e-11
.param cm4l1d=6.70e-05
.param cm4l1dsw=8.18e-11
.param cm4l1p1=1.06e-04
.param cm4l1p1sw=8.08e-11
.param cm5l1f=4.49e-05
.param cm5l1fsw=8.28e-11
.param cm5l1d=6.33e-05
.param cm5l1dsw=8.20e-11
.param cm5l1p1=1.02e-04
.param cm5l1p1sw=8.09e-11
.param crdll1f=3.97e-05
.param crdll1fsw=8.30e-11
.param crdll1d=5.80e-05
.param crdll1dsw=8.22e-11
.param crdll1p1=9.69e-05
.param crdll1p1sw=8.12e-11
.param cm2m1f=1.54e-04
.param cm2m1fsw=1.02e-10
.param cm2m1d=1.62e-04
.param cm2m1dsw=1.02e-10
.param cm2m1p1=1.73e-04
.param cm2m1p1sw=1.01e-10
.param cm2m1l1=2.42e-04
.param cm2m1l1sw=9.89e-11
.param cm3m1f=5.87e-05
.param cm3m1fsw=1.05e-10
.param cm3m1d=6.65e-05
.param cm3m1dsw=1.04e-10
.param cm3m1p1=7.78e-05
.param cm3m1p1sw=1.04e-10
.param cm3m1l1=1.47e-04
.param cm3m1l1sw=1.02e-10
.param cm4m1f=4.09e-05
.param cm4m1fsw=1.07e-10
.param cm4m1d=4.87e-05
.param cm4m1dsw=1.06e-10
.param cm4m1p1=6.00e-05
.param cm4m1p1sw=1.06e-10
.param cm4m1l1=1.29e-04
.param cm4m1l1sw=1.03e-10
.param cm5m1f=3.53e-05
.param cm5m1fsw=1.07e-10
.param cm5m1d=4.31e-05
.param cm5m1dsw=1.06e-10
.param cm5m1p1=5.44e-05
.param cm5m1p1sw=1.06e-10
.param cm5m1l1=1.23e-04
.param cm5m1l1sw=1.04e-10
.param crdlm1f=2.87e-05
.param crdlm1fsw=1.07e-10
.param crdlm1d=3.65e-05
.param crdlm1dsw=1.07e-10
.param crdlm1p1=4.78e-05
.param crdlm1p1sw=1.06e-10
.param crdlm1l1=1.17e-04
.param crdlm1l1sw=1.03e-10
.param cm3m2f=9.98e-05
.param cm3m2fsw=1.03e-10
.param cm3m2d=1.03e-04
.param cm3m2dsw=1.03e-10
.param cm3m2p1=1.07e-04
.param cm3m2p1sw=1.04e-10
.param cm3m2l1=1.19e-04
.param cm3m2l1sw=1.02e-10
.param cm3m2m1=2.10e-04
.param cm3m2m1sw=9.97e-11
.param cm4m2f=3.84e-05
.param cm4m2fsw=1.07e-10
.param cm4m2d=4.17e-05
.param cm4m2dsw=1.06e-10
.param cm4m2p1=4.56e-05
.param cm4m2p1sw=1.06e-10
.param cm4m2l1=5.79e-05
.param cm4m2l1sw=1.05e-10
.param cm4m2m1=1.49e-04
.param cm4m2m1sw=1.03e-10
.param cm5m2f=2.91e-05
.param cm5m2fsw=1.07e-10
.param cm5m2d=3.23e-05
.param cm5m2dsw=1.07e-10
.param cm5m2p1=3.62e-05
.param cm5m2p1sw=1.07e-10
.param cm5m2l1=4.85e-05
.param cm5m2l1sw=1.05e-10
.param cm5m2m1=1.39e-04
.param cm5m2m1sw=1.03e-10
.param crdlm2f=2.06e-05
.param crdlm2fsw=1.07e-10
.param crdlm2d=2.39e-05
.param crdlm2dsw=1.07e-10
.param crdlm2p1=2.78e-05
.param crdlm2p1sw=1.07e-10
.param crdlm2l1=4.01e-05
.param crdlm2l1sw=1.06e-10
.param crdlm2m1=1.31e-04
.param crdlm2m1sw=1.03e-10
.param cm4m3f=1.01e-04
.param cm4m3fsw=1.03e-10
.param cm4m3d=1.03e-04
.param cm4m3dsw=1.03e-10
.param cm4m3p1=1.04e-04
.param cm4m3p1sw=1.03e-10
.param cm4m3l1=1.09e-04
.param cm4m3l1sw=1.03e-10
.param cm4m3m1=1.21e-04
.param cm4m3m1sw=1.02e-10
.param cm4m3m2=1.71e-04
.param cm4m3m2sw=9.99e-11
.param cm5m3f=3.24e-05
.param cm5m3fsw=1.06e-10
.param cm5m3d=3.40e-05
.param cm5m3dsw=1.06e-10
.param cm5m3p1=3.57e-05
.param cm5m3p1sw=1.06e-10
.param cm5m3l1=4.00e-05
.param cm5m3l1sw=1.05e-10
.param cm5m3m1=5.27e-05
.param cm5m3m1sw=1.05e-10
.param cm5m3m2=1.02e-04
.param cm5m3m2sw=1.03e-10
.param crdlm3f=1.61e-05
.param crdlm3fsw=1.08e-10
.param crdlm3d=1.77e-05
.param crdlm3dsw=1.08e-10
.param crdlm3p1=1.94e-05
.param crdlm3p1sw=1.07e-10
.param crdlm3l1=2.37e-05
.param crdlm3l1sw=1.07e-10
.param crdlm3m1=3.64e-05
.param crdlm3m1sw=1.06e-10
.param crdlm3m2=8.57e-05
.param crdlm3m2sw=1.05e-10
.param cm5m4f=7.70e-05
.param cm5m4fsw=1.04e-10
.param cm5m4d=7.78e-05
.param cm5m4dsw=1.04e-10
.param cm5m4p1=7.85e-05
.param cm5m4p1sw=1.04e-10
.param cm5m4l1=8.01e-05
.param cm5m4l1sw=1.04e-10
.param cm5m4m1=8.35e-05
.param cm5m4m1sw=1.03e-10
.param cm5m4m2=8.92e-05
.param cm5m4m2sw=1.03e-10
.param cm5m4m3=1.57e-04
.param cm5m4m3sw=1.00e-10
.param crdlm4f=1.27e-05
.param crdlm4fsw=1.09e-10
.param crdlm4d=1.34e-05
.param crdlm4dsw=1.09e-10
.param crdlm4p1=1.41e-05
.param crdlm4p1sw=1.09e-10
.param crdlm4l1=1.57e-05
.param crdlm4l1sw=1.09e-10
.param crdlm4m1=1.91e-05
.param crdlm4m1sw=1.08e-10
.param crdlm4m2=2.49e-05
.param crdlm4m2sw=1.08e-10
.param crdlm4m3=9.25e-05
.param crdlm4m3sw=1.05e-10
.param crdlm5f=1.20e-05
.param crdlm5fsw=7.60e-11
.param crdlm5d=1.24e-05
.param crdlm5dsw=7.59e-11
.param crdlm5p1=1.27e-05
.param crdlm5p1sw=7.57e-11
.param crdlm5l1=1.35e-05
.param crdlm5l1sw=7.55e-11
.param crdlm5m1=1.50e-05
.param crdlm5m1sw=7.52e-11
.param crdlm5m2=1.70e-05
.param crdlm5m2sw=7.49e-11
.param crdlm5m3=2.53e-05
.param crdlm5m3sw=7.50e-11
.param crdlm5m4=7.39e-05
.param crdlm5m4sw=8.61e-11