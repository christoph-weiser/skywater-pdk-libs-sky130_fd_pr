* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b=-0.01
.param sky130_fd_pr__rf_pfet_01v8_b__toxe_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__overlap_mult=9.5435e-1
.param sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult=9.9626e-1
.param sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult=1.0009
.param sky130_fd_pr__rf_pfet_01v8_b__lint_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__wint_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__rshg_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__dlc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__xgw_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rd_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rs_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_0=-0.023953
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_0=-0.00025608
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_0='0.0054151+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_0=-1792.7
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_1=-0.0146
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_1=-0.00017534
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_1='-0.0013289+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_1=-3939.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_2=-0.017504
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_2=-0.00011528
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_2='0.0016874+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_2=-3705.2
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_3=-0.025672
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_3=-0.00043953
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_3='0.00554+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_3=-7604.3
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_4=-0.016429
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_4=-0.00040298
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_4='0.0090164+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_4=222.9
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_5=-0.018578
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_5=-0.00022966
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_5='0.0043185+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_5=12358.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_6=-0.026387
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_6=-0.00078906
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_6='0.013291+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_6=-3996.4
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_7=-0.00030611
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_7=-5407.7
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_7=-0.013695
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_7='0.0054619+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_8='0.0030552+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_8=-0.00032694
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_8=2232.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_8=-0.017831
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_0=-0.022271
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_0=-0.00043404
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_0='0.018047+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_0=-1656.1
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_1=-0.014049
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_1=-0.0002533
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_1='0.012426+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_1=876.35
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_2=-0.0001857
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_2='0.0094773+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_2=15921.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_2=-0.018595
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_3=-0.023461
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_3=-0.00053503
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_3='0.0064872+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_3=-2980.8
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_4=-0.00062465
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_4='0.022342+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_4=-1155.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_4=-0.012789
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_5='0.012097+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_5=-0.00033445
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_5=9117.5
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_5=-0.018599
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_6='0.017753+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_6=-0.00064602
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_6=-2850.2
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_6=-0.0251
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_7=-0.010953
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_7='0.0097164+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_7=-0.00057548
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_7=-3914.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_8=-0.016606
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_8='0.015491+sky130_fd_pr__pfet_01v8__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_8=-0.00044041
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_8=11410.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_8=0.0
.include "sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"