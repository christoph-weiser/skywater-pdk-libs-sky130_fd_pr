* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre=0.0
.subckt sky130_fd_pr__nfet_g5v0d10v5 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__nfet_g5v0d10v5 d g s b sky130_fd_pr__nfet_g5v0d10v5__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__nfet_g5v0d10v5__model.0 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.1 nmos lmin=8e-06 lmax=2.0e-05 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.2 nmos lmin=4e-06 lmax=8e-06 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.77946515163+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.78402092817277e-8 k1=0.88325 k2=-0.041896263236075 lk2=1.13681439985862e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=110499.05125 lvsat=-0.0380893386001013 ua=-1.0068597670945e-10 lua=3.35535078022468e-16 pua=1.50463276905253e-36 ub=1.5699538924075e-18 lub=7.88982559762499e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.040142764421725 lu0=9.36312121467687e-9 a0=1.03526353952745 la0=-7.40744697785784e-7 keta=-0.01724261541675 lketa=-3.20940767044453e-8 a1=0.0 a2=0.65972622 ags=0.144271878355825 lags=5.78097127669178e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0531863659525+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.22106050366323e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.2594415078275 lpclm=5.87261422536361e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=21.48369335 lbeta0=1.98064560720527e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414343723 lkt1=9.14144126402424e-8 kt2=-0.019151 at=237424.82 lat=-0.60942941760162 ute=-1.33731241 lute=3.0471470880081e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.3 nmos lmin=2e-06 lmax=4e-06 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.794841311733+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.16846121315708e-8 k1=0.88325 k2=-0.0431421107591 lk2=1.61911200094691e-08 wk2=2.11758236813575e-22 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=93689.627275 lvsat=0.0269839926783018 ua=1.084620204428e-10 lua=-4.74127223621206e-16 pua=5.64237288394698e-37 ub=1.534757614516e-18 lub=9.25235833783467e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.04229764858105 lu0=1.02104530684742e-9 a0=0.468487175688 la0=1.45338319974041e-6 keta=-0.0394484836965 lketa=5.38701910207224e-8 a1=0.0 a2=0.65972622 ags=0.120103548064 lags=1.51371143894173e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99177308345+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.84360433198061e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.603475506185 lpclm=-7.44577097299126e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=23.823078356 lbeta0=1.07501329220402e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=139879.712 lat=-0.231808796162592 ute=-1.22117518 lute=-1.4488049760162e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.4 nmos lmin=1e-06 lmax=2e-06 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.771193089784+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.25669103564979e-8 k1=0.88325 k2=-0.041376660105 lk2=1.28875363620403e-08 wk2=2.11758236813575e-22 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=120222.863623 lvsat=-0.0226660870387661 ua=-1.399951218104e-10 lua=-9.2040322941853e-18 ub=1.742611530568e-18 lub=5.36291064056405e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0415885387118 lu0=2.34796076769266e-9 a0=1.735670644457 la0=-9.17822461542362e-7 keta=0.003722446428 lketa=-2.69130234363772e-08 pketa=5.04870979341448e-29 a1=0.0 a2=0.65972622 ags=0.132297033427 lags=1.28554194150027e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.90313858535+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.85039263389194e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.09363295632 lpclm=2.09461185552807e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=27.013521388 lbeta0=4.78004511239749e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.38144241 lkt1=1.630301880081e-8 kt2=-0.019151 at=9030.072 lat=0.013042415040648 ute=-1.2986 ua1=3.0044e-9 ub1=-4.0140465482e-18 lub1=4.89416624400316e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.5 nmos lmin=8.0e-07 lmax=1e-06 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.778692706885+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=2.60329364538054e-8 k1=0.88325 k2=-0.0370474690875 lk2=9.11576765076259e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=64406.9201845 lvsat=0.025963051338536 ua=-1.687866137345e-10 lua=1.58802959212596e-17 ub=2.7598306144e-18 lub=-3.49951907760472e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.046078398434 lu0=-1.5637891065366e-9 a0=-0.794508418975001 la0=1.2865732758612e-6 keta=-0.08257223214 lketa=4.82704386138858e-8 a1=0.0 a2=0.65972622 ags=0.681252118 lags=-3.49717982688438e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.94838642105+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.79256959620228e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.99431721875 lpclm=2.02856898403097e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.757498935e-06 lalpha0=8.45931541737167e-12 alpha1=0.0 beta0=22.49179669 lbeta0=8.7195570600077e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.33588036 lkt1=-2.33925072032401e-8 kt2=-0.019151 at=7218.97499999999 lat=0.014620317002025 ute=-1.4714445575 lute=1.50589265120857e-7 ua1=6.3361047035e-09 lua1=-2.90271773758204e-15 ub1=-1.01824978865e-17 lub1=5.86362433683215e-24 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.6 nmos lmin=6e-07 lmax=8.0e-07 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.7620790286245+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.7184718463062e-8 k1=0.88325 k2=-0.0163350030855 lk2=-4.7872887408859e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90873.418244 lvsat=0.0081976527145792 ua=-3.0910151836e-10 lua=1.10065412816985e-16 ub=1.4358623288e-18 lub=5.38749888233959e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0392633339138 lu0=3.01076161706698e-9 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.93030213475+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.57867815417249e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.032041169 lpclm=-2.84684652072885e-9 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.667670055e-05 lalpha0=4.58658606117445e-13 alpha1=0.0 beta0=31.99952901 lbeta0=2.3375773097986e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.673 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210597e-8 ua1=2.0117e-9 ub1=-1.6826205e-18 lub1=1.581581400405e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.7 nmos lmin=5e-07 lmax=6e-07 wmin=2.0e-05 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.744876888751+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.52910720591901e-8 k1=0.88325 k2=-0.005538830514 lk2=-9.87488789965213e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=57681.402653 lvsat=0.0238390913336976 ua=2.31117104543e-10 lua=-1.44507751258448e-16 ub=-1.67464984888e-17 lub=9.1070237822806e-24 pub=2.24207754291971e-44 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0100033289894 lu0=1.67992755976462e-8 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.6229062217+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.90707759198702e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.0652282920000014 lpclm=4.52755020449628e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.946660103e-05 lalpha0=-5.56846688597823e-12 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960161999e-8 kt2=-0.019151 at=-3178.99199999997 lat=0.019593725769072 ute=-1.300956205 lute=8.74719900404651e-10 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=6.283858755e-18 lub1=-3.59597351056495e-24 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.8 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.9 nmos lmin=8e-06 lmax=2.0e-05 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.10 nmos lmin=4e-06 lmax=8e-06 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.77946515163+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.78402092817285e-8 k1=0.88325 k2=-0.041896263236075 lk2=1.13681439985862e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=110499.05125 lvsat=-0.0380893386001016 ua=-1.0068597670945e-10 lua=3.35535078022468e-16 ub=1.5699538924075e-18 lub=7.88982559762499e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.040142764421725 lu0=9.36312121467692e-9 a0=1.03526353952745 la0=-7.40744697785784e-7 keta=-0.01724261541675 lketa=-3.20940767044453e-8 a1=0.0 a2=0.65972622 ags=0.144271878355825 lags=5.78097127669174e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0531863659525+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.22106050366321e-07 wnfactor=-1.35525271560688e-20 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.2594415078275 lpclm=5.87261422536362e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=21.48369335 lbeta0=1.98064560720527e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414343723 lkt1=9.14144126402407e-8 kt2=-0.019151 at=237424.82 lat=-0.60942941760162 ute=-1.33731241 lute=3.04714708800811e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.11 nmos lmin=2e-06 lmax=4e-06 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.794841311733+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.16846121315712e-8 k1=0.88325 k2=-0.0431421107591 lk2=1.6191120009469e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=93689.627275 lvsat=0.0269839926783018 ua=1.084620204428e-10 lua=-4.74127223621206e-16 wua=-1.97215226305253e-31 pua=-3.76158192263132e-37 ub=1.534757614516e-18 lub=9.25235833783461e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.04229764858105 lu0=1.0210453068475e-9 a0=0.468487175688 la0=1.45338319974041e-6 keta=-0.0394484836965 lketa=5.38701910207224e-8 a1=0.0 a2=0.65972622 ags=0.120103548064 lags=1.51371143894173e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99177308345+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.84360433198062e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.603475506185 lpclm=-7.44577097299125e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=23.823078356 lbeta0=1.07501329220402e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=139879.712 lat=-0.231808796162592 ute=-1.22117518 lute=-1.44880497601619e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.12 nmos lmin=1e-06 lmax=2e-06 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.77367979289907+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=2.79136895327517e-08 wvth0=-4.95158988637212e-08 pvth0=9.26561801056196e-14 k1=0.88325 k2=-0.0413200142033192 lk2=1.27815382283332e-08 wk2=-1.12794837537031e-09 pk2=2.11066324587524e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=128018.171193753 lvsat=-0.0372529861727692 wvsat=-0.155222253491258 pvsat=2.90458244845238e-7 ua=-1.3837938841021e-10 lua=-1.22274588776902e-17 wua=-3.21729164811323e-17 pua=6.0203280409072e-23 ub=1.40172273049898e-18 lub=1.17417616318636e-24 wub=6.78786914517275e-24 pub=-1.27017390470822e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.041212726933814 lu0=3.05119517494302e-09 wu0=7.48326484081381e-09 pu0=-1.40029919839888e-14 a0=1.72726470445987 la0=-9.02092921976194e-07 wa0=1.67381330014738e-07 pa0=-3.1321080735811e-13 keta=0.003722446428 lketa=-2.69130234363771e-8 a1=0.0 a2=0.65972622 ags=0.14271676121324 lags=1.09056372307576e-07 wags=-2.07480412166652e-07 pags=3.88245853943136e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.896954308010535+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.93165302594317e-09 wnfactor=1.23142987769722e-07 pnfactor=-2.30430207577225e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.0936329563200002 lpclm=2.09461185552807e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=27.078482284423 lbeta0=4.65848761961412e-06 wbeta0=-1.29351877909377e-06 pbeta0=2.42048537371034e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.38144241 lkt1=1.63030188008102e-8 kt2=-0.019151 at=9030.072 lat=0.013042415040648 ute=-1.2986 ua1=3.0044e-9 ub1=-4.0140465482e-18 lub1=4.89416624400315e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.13 nmos lmin=8.0e-07 lmax=1e-06 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.766259191309647+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.43788218821206e-08 wvth0=2.47579494318565e-07 pvth0=-1.66185507345877e-13 k1=0.88325 k2=-0.037330698595904 lk2=9.30588290921323e-09 wk2=5.63974187684899e-09 pk2=-3.78562597715741e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=25430.3823307359 lvsat=0.0521257015840344 wvsat=0.776111267456294 pvsat=-5.20957703278628e-7 ua=-1.7686528073545e-10 lua=2.1303028437644e-17 wua=1.60864582405674e-16 pua=-1.07978903158564e-22 ub=4.46427461474509e-18 lub=-1.49404460299612e-24 wub=-3.39393457258637e-23 pub=2.27814803643745e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.04795745732393 lu0=-2.82509047487214e-09 wu0=-3.74163242040708e-08 pu0=2.51153708750643e-14 a0=-0.75247871898936 la0=1.25836121801314e-06 wa0=-8.36906650073692e-07 pa0=5.6176605670214e-13 keta=-0.08257223214 lketa=4.82704386138857e-8 a1=0.0 a2=0.65972622 ags=0.629153479068802 lags=-3.14747240193622e-07 wags=1.03740206083325e-06 pags=-6.96346796715769e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.97930780774732+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.86813984901172e-08 wnfactor=-6.15714938848662e-07 pnfactor=4.13293111267744e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.99431721875 lpclm=2.02856898403097e-06 ppclm=-1.29246970711411e-26 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.7574989349999e-06 lalpha0=8.4593154173717e-12 alpha1=0.0 beta0=22.1669922078853 lbeta0=8.9375791453868e-06 wbeta0=6.46759389546885e-06 pbeta0=-4.34131419398836e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.335880359999999 lkt1=-2.3392507203241e-8 kt2=-0.019151 at=7218.97499999992 lat=0.014620317002025 ute=-1.4714445575 lute=1.50589265120858e-7 ua1=6.3361047035e-09 lua1=-2.90271773758204e-15 ub1=-1.01824978865e-17 lub1=5.86362433683215e-24 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.14 nmos lmin=6e-07 lmax=8.0e-07 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.762079028624498+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.71847184630611e-8 k1=0.88325 k2=-0.0163350030855 lk2=-4.78728874088592e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90873.4182440001 lvsat=0.00819765271457917 ua=-3.0910151836e-10 lua=1.10065412816985e-16 ub=1.4358623288e-18 lub=5.3874988823396e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0392633339138 lu0=3.01076161706698e-9 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.930302134750002+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.57867815417249e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.032041169 lpclm=-2.84684652072885e-9 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.667670055e-05 lalpha0=4.58658606117452e-13 alpha1=0.0 beta0=31.99952901 lbeta0=2.33757730979859e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67299999995 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210601e-8 ua1=2.0117e-9 ub1=-1.6826205e-18 lub1=1.581581400405e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.15 nmos lmin=5e-07 lmax=6e-07 wmin=1.5e-05 wmax=2.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.743304651890174+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.60319745297211e-08 wvth0=3.13068017321588e-08 pvth0=-1.4753048555068e-14 k1=0.88325 k2=0.00339856099343888 lk2=-1.40865532110092e-08 wk2=-1.77963734917048e-07 pk2=8.38638084060446e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-82038.4154484896 lvsat=0.0896807981356617 wvsat=2.7821384629481 pvsat=-1.31105771141813e-6 ua=4.3450919388065e-10 lua=-2.40354442830011e-16 wua=-4.04999779197123e-15 pua=1.90852500948631e-21 ub=-5.20576097320163e-17 lub=2.57470671556451e-23 wub=7.03124310452735e-22 pub=-3.31341003182057e-28 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=-0.0269730246754204 lu0=3.42240494750097e-08 wu0=7.36283063836684e-07 pu0=-3.46966767285463e-13 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.420951289718227+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.94240220021891e-07 wnfactor=4.02138072954278e-06 pnfactor=-1.89503947637047e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-2.2111935290226 lpclm=1.52549831581014e-06 wpclm=4.53287213812499e-05 ppclm=-2.13607519924216e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.94666010299999e-05 lalpha0=-5.56846688597823e-12 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960161996e-8 kt2=-0.019151 at=-91047.1027569813 lat=0.0610007821503025 wat=1.74965337004669 pat=-8.24508403754172e-7 ute=-1.30095620499999 lute=8.74719900405922e-10 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=2.40862705578839e-18 lub1=-1.76980544939678e-24 wub1=7.71646521567969e-23 pub1=-3.63631478470211e-29 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.16 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.17 nmos lmin=8e-06 lmax=2.0e-05 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.18 nmos lmin=4e-06 lmax=8e-06 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.77946515163+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.78402092817285e-8 k1=0.88325 k2=-0.041896263236075 lk2=1.13681439985862e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=110499.05125 lvsat=-0.0380893386001011 ua=-1.0068597670945e-10 lua=3.35535078022468e-16 ub=1.5699538924075e-18 lub=7.88982559762499e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.040142764421725 lu0=9.36312121467671e-9 a0=1.03526353952745 la0=-7.40744697785788e-7 keta=-0.01724261541675 lketa=-3.20940767044453e-8 a1=0.0 a2=0.65972622 ags=0.144271878355825 lags=5.78097127669178e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0531863659525+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.22106050366321e-07 wnfactor=-6.7762635780344e-21 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.2594415078275 lpclm=5.87261422536359e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=21.48369335 lbeta0=1.98064560720526e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414343723 lkt1=9.14144126402424e-8 kt2=-0.019151 at=237424.82 lat=-0.60942941760162 ute=-1.33731241 lute=3.04714708800811e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.19 nmos lmin=2e-06 lmax=4e-06 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.794841311733+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.16846121315729e-8 k1=0.88325 k2=-0.0431421107591 lk2=1.61911200094691e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=93689.627275 lvsat=0.0269839926783018 ua=1.084620204428e-10 lua=-4.74127223621206e-16 pua=-5.64237288394698e-37 ub=1.534757614516e-18 lub=9.25235833783467e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.04229764858105 lu0=1.0210453068474e-9 a0=0.468487175687999 la0=1.45338319974041e-6 keta=-0.0394484836965 lketa=5.38701910207224e-8 a1=0.0 a2=0.65972622 ags=0.120103548064 lags=1.51371143894173e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99177308345+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.84360433198062e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.603475506185 lpclm=-7.44577097299125e-07 wpclm=3.3881317890172e-21 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=23.823078356 lbeta0=1.07501329220402e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=139879.712 lat=-0.231808796162592 ute=-1.22117518 lute=-1.4488049760162e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.20 nmos lmin=1e-06 lmax=2e-06 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.760206860778038+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=5.31247925078425e-08 wvth0=1.51396075670917e-07 pvth0=-2.83298544034532e-13 k1=0.88325 k2=-0.0388551222437599 lk2=8.16913133303554e-09 wk2=-3.78850778673631e-08 pk2=7.08921109936026e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=124903.084503763 lvsat=-0.031423908239906 wvsat=-0.108769245926898 pvsat=2.03533472517495e-7 ua=-1.36438597492065e-10 lua=-1.58591464161517e-17 wua=-6.11145107844858e-17 pua=1.14359978274872e-22 ub=1.47284195299952e-18 lub=1.04109495815523e-24 wub=5.72732023929309e-24 pub=-1.07171964518951e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0416193260451682 lu0=2.29035024721353e-09 wu0=1.41994992373892e-09 pu0=-2.65706851524715e-15 a0=2.70180785980979 la0=-2.72569803053634e-06 wa0=-1.43652673801289e-05 pa0=2.68808772976598e-11 keta=0.0322349791259957 lketa=-8.02668436347074e-08 wketa=-4.25186528951275e-07 pketa=7.95626465621313e-13 a1=0.0 a2=0.65972622 ags=0.0186394146530819 lags=3.41234990362153e-07 wags=1.6427942324673e-06 pags=-3.07406392235635e-12 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.873967183968361+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.60827959538607e-08 wnfactor=4.65933142035894e-07 pnfactor=-8.71873198636388e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.759362941970319 lpclm=-1.03628005852548e-06 wpclm=-9.92754396165371e-06 ppclm=1.85768272903489e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.24686355505463e-05 lalpha0=3.73942149076012e-12 walpha0=2.98001462319254e-11 palpha0=-5.57632554351745e-17 alpha1=0.0 beta0=27.4667189486524 lbeta0=3.93200325580486e-06 wbeta0=-7.0830079635085e-06 pbeta0=1.32540149046438e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.398714358569176 lkt1=4.86229971133435e-08 wkt1=2.5756392594577e-07 pkt1=-4.81964178350687e-13 kt2=-0.019151 at=9030.07200000001 lat=0.013042415040648 ute=-1.2986 ua1=3.0044e-9 ub1=-4.53255044424666e-18 lub1=1.45966237334257e-24 wub1=7.73206905689198e-24 pub1=-1.44685646340876e-29 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.21 nmos lmin=8.0e-07 lmax=1e-06 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.833623851914808+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.08391002671473e-08 wvth0=-7.56980378354606e-07 pvth0=5.08116266147124e-13 k1=0.88325 k2=-0.0496551583937005 lk2=1.75785656283459e-08 wk2=1.89425389336816e-07 pk2=-1.27150087763834e-13 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=41005.8157806848 lvsat=0.0416708320596573 wvsat=0.543846229634491 pvsat=-3.65051887026088e-7 ua=-1.86569235326177e-10 lua=2.78167206210788e-17 wua=3.05572553922429e-16 pua=-2.05112826667446e-22 ub=4.10867850224241e-18 lub=-1.2553539128437e-24 wub=-2.86366011964655e-23 pub=1.92220608237167e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0459244617671591 lu0=-1.46046050434972e-09 wu0=-7.09974961869419e-09 pu0=4.76564303380204e-15 a0=-5.62519449573898 la0=4.52912782871433e-06 wa0=7.18263369006448e-05 pa0=-4.82127822075257e-11 keta=-0.225134895629979 lketa=1.43964343417563e-07 wketa=2.12593264475638e-06 pketa=-1.42701315439892e-12 a1=0.0 a2=0.65972622 ags=1.24954021186959 lags=-7.31176251105557e-07 wags=-8.21397116233653e-06 pags=5.51355421697793e-12 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.09424342795819+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.55830899136088e-07 wnfactor=-2.32966571017948e-06 pnfactor=1.56376714096658e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-5.3229671470016 lpclm=4.2628952905205e-06 wpclm=4.96377198082686e-05 ppclm=-3.33188726818221e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.47493211822684e-05 lalpha0=1.75239466029304e-12 walpha0=-1.49000731159628e-10 palpha0=1.0001539978432e-16 alpha1=0.0 beta0=20.2258088867383 lbeta0=1.02405809790569e-05 wbeta0=3.54150398175429e-05 pbeta0=-2.37720267421673e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.249520617154119 lkt1=-8.13607073508517e-08 wkt1=-1.28781962972884e-06 pkt1=8.64437336078823e-13 kt2=-0.019151 at=7218.97500000003 lat=0.014620317002025 ute=-1.4714445575 lute=1.50589265120857e-7 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-7.58997840626669e-18 lub1=4.12341896840086e-24 wub1=-3.86603452844599e-23 pub1=2.59504088290862e-29 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.22 nmos lmin=6e-07 lmax=8.0e-07 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.762079028624499+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.71847184630628e-8 k1=0.88325 k2=-0.0163350030855 lk2=-4.78728874088589e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90873.4182440001 lvsat=0.00819765271457928 ua=-3.0910151836e-10 lua=1.10065412816985e-16 ub=1.4358623288e-18 lub=5.38749888233959e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0392633339138 lu0=3.01076161706698e-9 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.930302134749999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.5786781541724e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.032041169 lpclm=-2.84684652072885e-9 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.667670055e-05 lalpha0=4.58658606117439e-13 alpha1=0.0 beta0=31.99952901 lbeta0=2.33757730979859e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67300000001 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210601e-8 ua1=2.0117e-9 ub1=-1.6826205e-18 lub1=1.581581400405e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.23 nmos lmin=5e-07 lmax=6e-07 wmin=1.0e-05 wmax=1.5e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.764436184922886+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.60739297718538e-08 wvth0=-2.83812282102472e-07 pvth0=1.33743983630251e-13 k1=0.88325 k2=-0.0236368164258923 lk2=-1.34637492054614e-09 wk2=2.25195058641167e-07 pk2=-1.06121144629122e-13 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=109913.017988409 lvsat=-0.000774587308575936 wvsat=-0.0802927554470863 pvsat=3.78372383696406e-8 ua=6.00340129040334e-11 lua=-6.38863840714096e-17 wua=1.53427646610058e-15 pua=-7.23013976161705e-22 ub=-7.79113933186007e-18 lub=4.88689137780507e-24 wub=4.30108404315382e-23 pub=-2.02684714557985e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0148193505030347 lu0=1.45297688035394e-08 wu0=1.13063964819012e-07 pu0=-5.32803758452762e-14 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.811024954211717+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.04215162923149e-08 wnfactor=-1.79550229512622e-06 pnfactor=8.46114297057575e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=2.34165011302258 lpclm=-6.19988274910876e-07 wpclm=-2.25645031710239e-05 ppclm=1.06333190388165e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.946660103e-05 lalpha0=-5.56846688597823e-12 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960161998e-8 kt2=-0.019151 at=84689.1187569806 lat=-0.0218133306121583 wat=-0.870972262476876 pat=4.10437839941866e-7 ute=-1.300956205 lute=8.74719900405075e-10 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=7.583202255e-18 lub1=-4.20827744084845e-24 wub1=-2.35098870164458e-38 pub1=1.12103877145985e-44 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.24 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.25 nmos lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.785543+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.040452 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=105660.0 ua=-5.8058e-11 ub=1.67019e-18 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0413323 a0=0.9411558 keta=-0.02132 a1=0.0 a2=0.65972622 ags=0.1516163 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99956+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.33405 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=24.0 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=160000.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.26 nmos lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.779465151629999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.78402092817285e-8 k1=0.88325 k2=-0.041896263236075 lk2=1.13681439985864e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=110499.05125 lvsat=-0.0380893386001011 ua=-1.0068597670945e-10 lua=3.35535078022468e-16 ub=1.5699538924075e-18 lub=7.88982559762493e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.040142764421725 lu0=9.36312121467692e-9 a0=1.03526353952745 la0=-7.40744697785781e-7 keta=-0.01724261541675 lketa=-3.20940767044453e-8 a1=0.0 a2=0.65972622 ags=0.144271878355825 lags=5.78097127669182e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0531863659525+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.22106050366321e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.2594415078275 lpclm=5.8726142253636e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=21.48369335 lbeta0=1.98064560720528e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414343723 lkt1=9.14144126402424e-8 kt2=-0.019151 at=237424.82 lat=-0.60942941760162 ute=-1.33731241 lute=3.04714708800811e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.27 nmos lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.794841311733+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.16846121315712e-8 k1=0.88325 k2=-0.0431421107591 lk2=1.61911200094691e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=93689.627275 lvsat=0.0269839926783018 ua=1.084620204428e-10 lua=-4.74127223621205e-16 wua=-1.97215226305253e-31 pua=-7.52316384526264e-37 ub=1.534757614516e-18 lub=9.25235833783464e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.04229764858105 lu0=1.0210453068475e-09 wu0=2.11758236813575e-22 a0=0.468487175688 la0=1.45338319974041e-6 keta=-0.0394484836965 lketa=5.38701910207224e-8 a1=0.0 a2=0.65972622 ags=0.120103548064 lags=1.51371143894172e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.99177308345+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.84360433198062e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.603475506185 lpclm=-7.44577097299125e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=23.823078356 lbeta0=1.07501329220401e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=139879.712 lat=-0.231808796162592 ute=-1.22117518 lute=-1.44880497601619e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.28 nmos lmin=1e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.775480466745001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=2.45441948046198e-8 k1=0.88325 k2=-0.0426771615457 lk2=1.53210879784372e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=113929.88988 lvsat=-0.0108904165589411 ua=-1.42604140109e-10 lua=-4.32193028409483e-18 ub=2.050643142323e-18 lub=-4.01103171556335e-26 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.04176257781396 lu0=2.02229166412768e-9 a0=1.252566638716 la0=-1.38184387355667e-8 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.184372850479 lags=3.11077901738257e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.920972888620001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.18762058241777e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.24217817472 lpclm=8.37844742211227e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.5475025837e-05 lalpha0=-1.88625927525372e-12 alpha1=0.0 beta0=26.752149088 lbeta0=5.26913567642178e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=9030.072 lat=0.013042415040648 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.29 nmos lmin=8.0e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.757255822080001+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.04222524471981e-8 k1=0.88325 k2=-0.030544961884 lk2=4.75101821297807e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=95871.7888995002 lvsat=0.0048425413974108 ua=-1.557415222415e-10 lua=7.12389566240659e-18 ub=1.219672555625e-18 lub=6.83865327769718e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0452082029231999 lu0=-9.79678201671659e-10 a0=1.62101160973 la0=-3.34822803726776e-7 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.42087303274 lags=-1.7494086511943e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.859214904699998+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.92988184426676e-9 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.315261563550001 lpclm=9.01517986978867e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-2.82630250000052e-07 lalpha0=1.18424567716403e-11 alpha1=0.0 beta0=23.79865819 lbeta0=7.84233803988621e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.379442410000001 lkt1=5.84812680080982e-9 kt2=-0.019151 at=7218.97500000003 lat=0.014620317002025 ute=-1.4714445575 lute=1.50589265120858e-7 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-1.14902306275e-17 lub1=6.74142816963373e-24 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.30 nmos lmin=6e-07 lmax=8.0e-07 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.7620790286245+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.7184718463062e-8 k1=0.88325 k2=-0.0163350030855 lk2=-4.78728874088589e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90873.4182440001 lvsat=0.00819765271457917 ua=-3.0910151836e-10 lua=1.10065412816985e-16 ub=1.4358623288e-18 lub=5.3874988823396e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0392633339138 lu0=3.01076161706698e-9 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.930302134750001+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.57867815417257e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.032041169 lpclm=-2.8468465207297e-9 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.667670055e-05 lalpha0=4.58658606117452e-13 alpha1=0.0 beta0=31.9995290100001 lbeta0=2.33757730979859e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67299999995 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210601e-8 ua1=2.0117e-9 ub1=-1.6826205e-18 lub1=1.581581400405e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.31 nmos lmin=5e-07 lmax=6e-07 wmin=7e-06 wmax=1.0e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.573471179287965+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.26064469992261e-07 wvth0=1.60908403237241e-06 pvth0=-7.58266368499211e-13 k1=0.88325 k2=0.0188693365944579 lk2=-2.1377016976009e-08 wk2=-1.96137321745554e-07 pk2=9.24279476366968e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=95292.1725078621 lvsat=0.00611535453652268 wvsat=0.0646329833426869 pvsat=-3.0457711703391e-8 ua=2.89790451857094e-10 lua=-1.72157038120089e-16 wua=-7.43130931527799e-16 pua=3.50193763304092e-22 ub=-9.91432573282076e-18 lub=5.8874238605802e-24 wub=6.40564330518161e-23 pub=-3.01860175677709e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0131249340971502 lu0=1.53282472850649e-08 wu0=1.29859474337739e-07 pu0=-6.11951085463907e-14 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.426050302860896+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.91837355969529e-07 wnfactor=2.02046962226973e-06 pnfactor=-9.52128125268e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.065228292000004 lpclm=4.52755020449628e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.946660103e-05 lalpha0=-5.56846688597823e-12 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960162005e-8 kt2=-0.019151 at=-85294.7451068157 lat=0.058290035378881 wat=0.813953351816592 pat=-3.83568191463403e-7 ute=-1.300956205 lute=8.74719900404228e-10 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=9.29394711139199e-18 lub1=-5.01445055771948e-24 wub1=-1.6957361496179e-23 pub1=7.99100398882087e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.32 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.771719877848+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=9.55491249113593e-8 k1=0.88325 k2=-0.04029235129 wk2=-1.10353466937412e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=119095.05298 wvsat=-0.0928666867919588 ua=-3.738485518748e-10 wua=2.18282892642652e-15 ub=2.08395033364e-18 wub=-2.8600223138891e-24 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0403933199718 wu0=6.49048160156592e-9 a0=1.225977695109 wa0=-1.9687652712613e-6 keta=-0.017068432046 wketa=-2.93879771182598e-8 a1=0.0 a2=0.65972622 ags=0.1665675244982 wags=-1.03346870659724e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.9517881937+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=3.30211527989689e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.6505228659 wpclm=-2.18754526382886e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.3704519974e-05 walpha0=-6.3852213715641e-11 alpha1=0.0 beta0=26.66490539 wbeta0=-1.84205402503245e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=179649.072 wat=-0.135819651615296 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.33 nmos lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.771719877848+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=9.55491249113593e-8 k1=0.88325 k2=-0.04029235129 wk2=-1.10353466937434e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=119095.05298 wvsat=-0.0928666867919588 ua=-3.738485518748e-10 wua=2.18282892642652e-15 ub=2.08395033364e-18 wub=-2.86002231388909e-24 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0403933199718 wu0=6.49048160156571e-9 a0=1.225977695109 wa0=-1.9687652712613e-6 keta=-0.017068432046 wketa=-2.93879771182597e-8 a1=0.0 a2=0.65972622 ags=0.1665675244982 wags=-1.03346870659724e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.9517881937+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=3.30211527989686e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.6505228659 wpclm=-2.18754526382886e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.3704519974e-05 walpha0=-6.3852213715641e-11 alpha1=0.0 beta0=26.66490539 wbeta0=-1.84205402503245e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=179649.072 wat=-0.135819651615296 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.34 nmos lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.757864251004603+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.09060978090448e-07 wvth0=1.49311214164111e-07 pvth0=-4.23174361171891e-13 k1=0.88325 k2=-0.0435843123278388 lk2=2.59118186914395e-08 wk2=1.1668247719428e-08 pk2=-1.00529777181817e-13 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=142071.161000176 lvsat=-0.180850483468836 wvsat=-0.218234883918629 pvsat=9.86803293319524e-7 ua=-5.22074609204903e-10 lua=1.16672301972506e-15 wua=2.91275115996208e-15 pua=-5.74539381141667e-21 ub=2.10107025393002e-18 lub=-1.34755018503489e-25 wub=-3.6712186300285e-24 pub=6.38512170264544e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0385550815373545 lu0=1.44692177329832e-08 wu0=1.09744895957817e-08 pu0=-3.52947075683999e-14 a0=1.53821622703315 la0=-2.45770473426116e-06 wa0=-3.47654376735963e-06 pa0=1.18680879174075e-11 keta=-0.00297644455675386 lketa=-1.10921429696841e-07 wketa=-9.8611596318084e-08 pketa=5.44875789614044e-13 a1=0.0 a2=0.65972622 ags=0.187156785058922 lags=-1.62063031885241e-07 wags=-2.96431968286806e-07 pags=1.51981933693129e-12 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.962793664778417+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-8.66267151767493e-08 wnfactor=6.24818575759177e-07 pnfactor=-2.31892307329213e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.392665919413889 lpclm=2.02965416931628e-06 wpclm=-9.20882837027425e-07 ppclm=-9.97020522699896e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=3.53949584007005e-05 lalpha0=-9.20182582522203e-11 walpha0=-1.44659657158493e-10 palpha0=6.36054861932559e-16 alpha1=0.0 beta0=26.7538692799886 lbeta0=-7.00256218397481e-07 wbeta0=-3.64288684352302e-05 pbeta0=1.41747891150485e-10 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414343723 lkt1=9.14144126402441e-8 kt2=-0.019151 at=276090.465284588 lat=-0.759113448918774 wat=-0.267267302600009 pat=1.03465613978456e-6 ute=-1.33731241 lute=3.04714708800805e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.35 nmos lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.796383011754139+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-4.00544277923458e-08 wvth0=-1.0656643721712e-08 pvth0=1.9609976895787e-13 k1=0.88325 k2=-0.0404004519616682 lk2=1.35863279036445e-08 wk2=-1.89510803724064e-08 pk2=1.80050211197436e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=72941.7551968921 lvsat=0.086766106582473 wvsat=0.143414852233598 pvsat=-4.13229992912158e-7 ua=1.24566203184841e-10 lua=-1.33657940547143e-15 wua=-1.11316427033966e-16 pua=5.96150061813349e-21 ub=1.29244290326546e-18 lub=2.99563633511051e-24 wub=1.67494422450636e-24 pub=-1.43111631325069e-29 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0431899018304934 lu0=-3.47328861344819e-09 wu0=-6.16749358402389e-09 pu0=3.10660405385748e-14 a0=0.271915731940941 la0=2.4444496606601e-06 wa0=1.3587545003266e-06 pa0=-6.85051698368839e-12 keta=-0.0512482674195869 lketa=7.59504301144952e-08 wketa=8.15632674360142e-08 pketa=-1.52624530120235e-13 a1=0.0 a2=0.65972622 ags=0.100322889281791 lags=1.74091905636918e-07 wags=1.36729214719185e-07 pags=-1.57051994330005e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.01933864672402+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.05525967628839e-07 wnfactor=-1.90540560921e-07 pnfactor=8.37528646348754e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.58169351829319 lpclm=-2.57335822159682e-06 wpclm=-6.76170506211904e-06 ppclm=1.26410252444869e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=8.96645617743293e-06 lalpha0=1.02928431230843e-11 walpha0=3.80212330473281e-11 palpha0=-7.11468901487154e-17 alpha1=0.0 beta0=23.7707827794674 lbeta0=1.08479905489666e-05 wbeta0=3.6148104020793e-07 pbeta0=-6.76418143159869e-13 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207284e-8 kt2=-0.019151 at=149071.749284588 lat=-0.267393387772218 wat=-0.0635378251770646 pat=2.45970233876284e-7 ute=-1.22117518 lute=-1.44880497601622e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.36 nmos lmin=1e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.76674014069943+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.54145278829376e-08 wvth0=6.04154760343575e-08 pvth0=6.31067045134022e-14 k1=0.88325 k2=-0.0418321007113529 lk2=1.62652877416533e-08 wk2=-5.84128696331073e-09 pk2=-6.52656180888616e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=125851.002044453 lvsat=-0.0122398453978039 wvsat=-0.0824019221387595 pvsat=9.32761378114751e-9 ua=-9.80164489100602e-10 lua=7.30637959891474e-16 wua=5.78944159840348e-15 pua=-5.0802397301441e-21 ub=3.5975866961358e-18 lub=-1.31784324100398e-24 wub=-1.06928884248265e-23 pub=8.83203240206339e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0378687997879624 lu0=6.48377569371948e-09 wu0=2.69148372482059e-08 pu0=-3.08389732902586e-14 a0=1.56496519129665 la0=2.48424972858563e-08 wa0=-2.15938251824955e-06 pa0=-2.6723475091093e-13 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.227297607951765 lags=-6.35083939018029e-08 wags=-2.96707427486753e-07 pags=6.54012421468075e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.892539148046982+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.82535469249148e-08 wnfactor=1.96541635083172e-07 pnfactor=1.13204570815709e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.144423402787071 lpclm=1.16120546612968e-07 wpclm=-2.67229371295164e-06 ppclm=4.98875106205959e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.89085834882014e-05 lalpha0=-6.44485031280456e-11 walpha0=-2.31101710678555e-10 palpha0=4.3244699619185e-16 alpha1=0.0 beta0=32.7438260864232 lbeta0=-5.94273598178465e-06 wbeta0=-4.14160771825367e-05 pbeta0=7.74994616831273e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=3485.30528458799 lat=0.00503393528478628 wat=0.0383269135344075 pat=5.53567583450909e-8 ute=-1.2986 ua1=3.0044e-9 ub1=-3.1105346073118e-18 lub1=-1.20127196337926e-24 wub1=-4.43743684098607e-24 pub1=8.30351375176364e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.37 nmos lmin=8.0e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.702944891356772+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=7.09955647154831e-08 wvth0=3.75411708488389e-07 pvth0=-2.11330928046077e-13 k1=0.88325 k2=-0.0238655522812298 lk2=6.1209412084442e-10 wk2=-4.61698692561207e-08 pk2=2.86093525564839e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=177193.208695701 lvsat=-0.0569712808628438 wvsat=-0.562115447771848 pvsat=4.27273705567245e-7 ua=-1.15877413166261e-10 lua=-2.23643764326361e-17 wua=-2.75551405509285e-16 pua=2.03830839577856e-22 ub=1.56692602899635e-18 lub=4.51351589295268e-25 wub=-2.40030907187358e-24 pub=1.6071972740173e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0452377602845098 lu0=6.36351817471374e-11 wu0=-2.04308402745504e-10 pu0=-7.21166171417769e-15 a0=3.17518842658171 la0=-1.37805000444714e-06 wa0=-1.0742886677466e-05 pa0=7.21106599626893e-12 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.134781155488503 lags=1.70957326587422e-08 wags=1.97754372818545e-06 pags=-1.32740842965093e-12 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.822947022531256+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.62203389846513e-09 wnfactor=2.5069332134278e-07 pnfactor=6.60254015272008e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-3.89163954168359 lpclm=3.63250406241653e-06 wpclm=2.47208830541575e-05 ppclm=-1.88773076576934e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-0.000143594339528013 lalpha0=1.03267936023524e-10 walpha0=9.90608942067715e-10 palpha0=-6.31957414617463e-16 alpha1=0.0 beta0=-6.15972680211615 lbeta0=2.79516343403792e-05 wbeta0=0.000207080385912684 pbeta0=-1.39000845320416e-10 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.379442409999999 lkt1=5.84812680080982e-9 kt2=-0.019151 at=-56977.5642688201 lat=0.0577116662173671 wat=0.443743684098609 pat=-2.97858954258034e-7 ute=-1.4714445575 lute=1.50589265120857e-7 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-1.31338326407617e-17 lub1=7.53143623858166e-24 wub1=1.13610176010044e-23 pub1=-5.46074749473064e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.38 nmos lmin=6e-07 lmax=8.0e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.732666972717976+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=5.10448851005082e-08 wvth0=2.03304012856886e-07 pvth0=-9.58051863226916e-14 k1=0.88325 k2=-0.0146121556403028 lk2=-5.59916509380809e-09 wk2=-1.19087832643186e-08 pk2=5.61190693426083e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=54735.6626698368 lvsat=0.0252272447891035 wvsat=0.249793851447111 pvsat=-1.17713104349788e-7 ua=-3.22750756636352e-10 lua=1.16497493511571e-16 wua=9.43471929620032e-17 pua=-4.44602655586075e-23 ub=1.43874748002401e-18 lub=5.37390286686004e-25 wub=-1.9942938480902e-26 pub=9.39793027267578e-33 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0445791013947086 lu0=5.05754033596132e-10 wu0=-3.67440094537249e-08 pu0=1.73152837589829e-14 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.760820108562177+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.40800979610499e-08 wnfactor=1.17150518619325e-06 pnfactor=-5.52061275446896e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=2.68391389408647 lpclm=-7.81277001363203e-07 wpclm=-1.1418186977688e-05 ppclm=5.38071784955268e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-7.17937842799416e-06 lalpha0=1.17006211197864e-11 walpha0=1.64899611325062e-10 palpha0=-7.77074577404335e-17 alpha1=0.0 beta0=31.99952901 lbeta0=2.33757730979856e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67300000001 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210592e-8 ua1=2.0117e-9 ub1=-3.2488454501793e-18 lub1=8.96227551787944e-25 wub1=1.0826166603926e-23 pub1=-5.10173357660068e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.39 nmos lmin=5e-07 lmax=6e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.821311984965273+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=9.2717208840796e-09 wvth0=-1.04058037805055e-07 pvth0=4.90364137932968e-14 k1=0.88325 k2=0.0108105705932454 lk2=-1.75793960268315e-08 wk2=-1.40432971395884e-07 pk2=6.61777738735678e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=115704.818307311 lvsat=-0.00350392108265551 wvsat=-0.076464695012179 pvsat=3.60332993422343e-8 ua=1.86475825870552e-10 lua=-1.23470950455565e-16 wua=-2.89925483890538e-17 pua=1.36624774954067e-23 ub=-1.01016470443302e-18 lub=1.69141811340172e-24 wub=2.50848570844438e-24 pub=-1.18210131373303e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0286921172684598 lu0=7.99235232023363e-09 wu0=2.22549322525553e-08 pu0=-1.04874365296263e-14 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.231988752400378+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.83287115070092e-07 wnfactor=3.36187506754833e-06 pnfactor=-1.58425336870654e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.0652282919999969 lpclm=4.52755020449628e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.94666010299999e-05 lalpha0=-5.56846688597823e-12 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960162e-8 kt2=-0.019151 at=119994.637660224 lat=-0.0384507386456416 wat=-0.605061879423769 pat=2.85129965121537e-7 ute=-1.300956205 lute=8.74719900405922e-10 ua1=-1.67360940700001e-09 lua1=1.73666889026409e-15 ub1=6.84072025500001e-18 lub1=-3.85838948068646e-24 pub1=5.60519385729927e-45 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.40 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.788903799362+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=1.11370971436263e-8 k1=0.88325 k2=-0.042712850072 wk2=1.07866040414833e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=132466.666244 wvsat=-0.158551634737081 ua=3.864226169134e-10 wua=-1.55182680733435e-15 ub=1.09854105674e-18 wub=1.98057214392992e-24 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0444767405846 wu0=-1.35683748052319e-8 a0=0.6282718728966 wa0=9.67325912606365e-7 keta=-0.012451800614 wketa=-5.20661079694674e-8 a1=0.0 a2=0.65972622 ags=0.1103186605862 wags=1.72962623571549e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0266547035+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=-3.75528323725381e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.80558997744 wpclm=4.96527126089923e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=5.229480026e-06 walpha0=2.6902133819641e-11 alpha1=0.0 beta0=21.62632141 wbeta0=6.33033459994216e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=207915.5456 wat=-0.274672145353421 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.41 nmos lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.788903799362+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=1.11370971436288e-8 k1=0.88325 k2=-0.042712850072 wk2=1.07866040414833e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=132466.666244 wvsat=-0.158551634737081 ua=3.864226169134e-10 wua=-1.55182680733435e-15 ub=1.09854105674e-18 wub=1.98057214392991e-24 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0444767405846 wu0=-1.35683748052319e-8 a0=0.6282718728966 wa0=9.67325912606365e-7 keta=-0.012451800614 wketa=-5.20661079694674e-8 a1=0.0 a2=0.65972622 ags=0.1103186605862 wags=1.72962623571548e-7 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0266547035+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=-3.75528323725381e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.80558997744 wpclm=4.96527126089923e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=5.229480026e-06 walpha0=2.6902133819641e-11 alpha1=0.0 beta0=21.62632141 wbeta0=6.33033459994213e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.40273 kt2=-0.019151 at=207915.5456 wat=-0.274672145353421 ute=-1.2986 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.42 nmos lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.787545632204452+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.06904610153446e-08 wvth0=3.50831510028937e-09 pvth0=6.00479819995801e-14 k1=0.88325 k2=-0.0425014978365724 lk2=-1.66360438093944e-09 wk2=6.3491727440436e-09 pk2=3.492809116309e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=137534.155426418 lvsat=-0.0398874286197057 wvsat=-0.195947896622837 pvsat=2.94354989801892e-7 ua=3.88072374623164e-10 lua=-1.29856405251651e-17 wua=-1.55813474399305e-15 pua=4.9651289653366e-23 ub=9.50171841752357e-19 lub=1.16784984814856e-24 wub=1.98230281136262e-24 pub=-1.36225004536179e-32 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0429818378875372 lu0=1.1766739400131e-08 wu0=-1.07709239670175e-08 pu0=-2.20194097332372e-14 a0=0.634514180365996 la0=-4.91347064877203e-08 wa0=9.6268287801792e-07 pa0=3.65464442169823e-14 keta=-0.012451800614 wketa=-5.20661079694674e-8 a1=0.0 a2=0.65972622 ags=0.100859071335681 lags=7.44587067518483e-08 wags=1.27485529309037e-07 pags=3.57961168919949e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.10903483204654+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.48433845400792e-07 wnfactor=-9.35572304946693e-08 pnfactor=4.40824114679245e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.80558997744 wpclm=4.96527126089923e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-7.27692075742253e-06 lalpha0=9.84408946089076e-11 walpha0=6.49560493298215e-11 palpha0=-2.99531539974269e-16 alpha1=0.0 beta0=16.9275226431835 lbeta0=3.69853775041156e-05 wbeta0=1.1840779705655e-05 pbeta0=-4.33740414443368e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414343723 lkt1=9.14144126402433e-8 kt2=-0.019151 at=303528.293554552 lat=-0.752590981822539 wat=-0.40204926840005 pat=1.00261603338667e-6 ute=-1.33731241 lute=3.04714708800811e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.43 nmos lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.795809023991763+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-2.12991200707547e-08 wvth0=-7.83706200420227e-09 pvth0=1.03968671006953e-13 k1=0.88325 k2=-0.0476736940599409 lk2=1.83592136990097e-08 wk2=1.67770340431912e-08 pk2=-5.44067304048325e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=144686.472175751 lvsat=-0.0675757704647103 wvsat=-0.209014425150707 pvsat=3.44938670766656e-7 ua=4.60533054954615e-10 lua=-2.93498397112168e-16 wua=-1.76167564204337e-15 pua=8.37607159362556e-22 ub=1.14924415198795e-18 lub=3.97192958799783e-25 wub=2.3783748680468e-24 pub=-1.54691288524377e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0456765152334241 lu0=1.33499397696265e-09 wu0=-1.83824050316114e-08 pu0=7.44646783474193e-15 a0=0.169965732125598 la0=1.74924429282689e-06 wa0=1.85956022201951e-06 pa0=-3.43548190185309e-12 keta=-0.0409264341123324 lketa=1.10232168658718e-07 wketa=3.08596559794542e-08 pketa=-3.21025617355388e-13 a1=0.0 a2=0.65972622 ags=0.0299671861991108 lags=3.48898279059828e-07 wags=4.82335283589735e-07 pags=-1.01574774869142e-12 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.00490206193018+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.45310796282782e-07 wnfactor=-1.1962418740894e-07 pnfactor=5.41735587031003e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.80558997744 wpclm=4.96527126089923e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.15994685360112e-05 lalpha0=-1.33465675557941e-11 walpha0=-2.40355093053205e-11 palpha0=4.49762304679972e-17 alpha1=0.0 beta0=24.0458347390387 lbeta0=9.42867586784484e-06 wbeta0=-9.89647899131657e-07 pbeta0=6.29563594684507e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207288e-8 kt2=-0.019151 at=178883.79821147 lat=-0.270062101026089 wat=-0.209982599135021 pat=2.59079668594454e-7 ute=-1.22117518 lute=-1.4488049760162e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.44 nmos lmin=1e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.767389029662501+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.18815385379254e-08 wvth0=5.72279595455082e-08 pvth0=-1.77836649827536e-14 k1=0.88325 k2=-0.0473971059689752 lk2=1.7841650723083e-08 wk2=2.1495510283539e-08 pk2=-1.42700792389479e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123415.594228365 lvsat=-0.0277728315435654 wvsat=-0.0704385462568395 pvsat=8.56298045694158e-8 ua=7.0388624735592e-10 lua=-7.48870868214379e-16 wua=-2.48306694466832e-15 pua=2.18750414187778e-21 ub=7.56586994595272e-19 lub=1.13194913065643e-24 wub=3.26286349706058e-24 pub=-3.20200427188815e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0470268366949977 lu0=-1.19178290511392e-09 wu0=-1.80718943930424e-08 pu0=6.86542759691559e-15 a0=1.12515210048107 la0=-3.81396022809769e-08 wa0=1.09725374491038e-09 pa0=4.21502013640429e-14 keta=0.042936376223923 lketa=-4.66953604177069e-08 wketa=-2.63279763840738e-07 pketa=2.29380124728368e-13 a1=0.0 a2=0.65972622 ags=0.171123031418018 lags=8.47616740965546e-08 wags=-2.07628527664786e-08 pags=-7.43298889180789e-14 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.888755977586946+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.79734812702567e-08 wnfactor=2.15125582272553e-07 pnfactor=-8.46619067375679e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-2.2910123007348 lpclm=2.77958315366449e-06 wpclm=9.29121915951634e-06 ppclm=-8.09489107175618e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-1.09847977125113e-05 lalpha0=4.76264474033574e-11 walpha0=6.3110629205508e-11 palpha0=-1.18095196905144e-16 alpha1=0.0 beta0=21.3820242140149 lbeta0=1.4413307338501e-05 wbeta0=1.43961385776347e-05 pbeta0=-2.24948785257255e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=30923.504569176 lat=0.00680726680941053 wat=-0.096456874788897 pat=4.66456786432879e-8 ute=-1.2986 ua1=3.0044e-9 ub1=-4.0138723e-18 lub1=4.89090564024298e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.45 nmos lmin=8.0e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.746719642630565+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=4.98895559650175e-08 wvth0=1.6037839859818e-07 pvth0=-1.07652556653441e-13 k1=0.88325 k2=-0.0378017468121645 lk2=9.48178041594411e-09 wk2=2.22884531799643e-08 pk2=-1.49609236009724e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=38068.1195877474 lvsat=0.046585387609801 wvsat=0.121304275450302 pvsat=-8.14244031575366e-8 ua=-1.96557757805301e-10 lua=3.56328672862879e-17 wua=1.20772069690043e-16 pua=-8.10671648308141e-23 ub=1.44397060542303e-18 lub=5.33072346175241e-25 wub=-1.79631907922797e-24 pub=1.20576301506006e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0542343032921631 lu0=-7.47122331069485e-09 wu0=-4.4397738729865e-08 pu0=2.98015825427732e-14 a0=0.944361943471263 la0=1.19372194902406e-07 wa0=2.15530869070061e-07 pa0=-1.44673156085455e-13 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.631423524311101 lags=-3.16270987632107e-07 wags=-4.62096687625992e-07 pags=3.10178242698758e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.76938148374286+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.60304721209582e-08 wnfactor=5.13821603435778e-07 pnfactor=-3.44898126911836e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.14083894975 lpclm=-2.1038636165914e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=0.000122303630227557 lalpha0=-6.84998958435754e-11 walpha0=-3.1555314602754e-10 palpha0=2.11812209292672e-16 alpha1=0.0 beta0=46.1261516737177 lbeta0=-7.14479101361789e-06 wbeta0=-4.97618617760424e-05 pbeta0=3.34022018604125e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37944241 lkt1=5.84812680080982e-9 kt2=-0.019151 at=71415.5142688201 lat=-0.028471032213317 wat=-0.186957527023328 pat=1.25493557396666e-7 ute=-1.4714445575 lute=1.50589265120858e-7 ua1=6.3361047035e-09 lua1=-2.90271773758204e-15 ub1=-1.08210480775e-17 lub1=6.41978119558918e-24 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.46 nmos lmin=6e-07 lmax=8.0e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.802512670783581+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.24389879545584e-08 wvth0=-1.3979677468845e-07 pvth0=9.38373268386504e-14 k1=0.88325 k2=-0.00975391501163381 lk2=-9.34507424967596e-09 wk2=-3.57737632408292e-08 pk2=2.40128166115374e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=102261.751493564 lvsat=0.00349598993570832 wvsat=0.0163329661531555 pvsat=-1.09633565336103e-8 ua=-5.31735783400807e-10 lua=2.60618100365041e-16 wua=1.12093765241618e-15 pua=-7.52419310745486e-22 ub=1.0782805490825e-18 lub=7.78538505283317e-25 wub=1.75076723144131e-24 pub=-1.17518674719989e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0312009256346633 lu0=7.98972414150303e-09 wu0=2.89731752307217e-08 pu0=-1.94479831150449e-14 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.04541768039216+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.09256340554111e-07 wnfactor=-2.26514358784861e-07 pnfactor=1.52045724705108e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.24742116377844 lpclm=-2.81928713585801e-07 wpclm=-4.36174970636323e-06 ppclm=2.92778523464896e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.83726470422297e-05 lalpha0=-5.44956875927327e-12 walpha0=-9.74146572750361e-12 palpha0=6.53887119639528e-18 alpha1=0.0 beta0=31.99952901 lbeta0=2.33757730979859e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67300000004 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210601e-8 ua1=2.0117e-9 ub1=-1.61447928510402e-18 lub1=2.39954752812507e-25 wub1=2.79772199094395e-24 pub1=-1.87794570692321e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.47 nmos lmin=5e-07 lmax=6e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.812107774403211+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=7.9173817297407e-09 wvth0=-5.88444887957754e-08 pvth0=5.56892906823021e-14 k1=0.88325 k2=-0.0413202322426017 lk2=5.5302686485626e-09 wk2=1.15647503188956e-07 pk2=-4.73430924021011e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=125465.541550129 lvsat=-0.00743858729433722 wvsat=-0.12441198345473 pvsat=5.53614342645595e-8 ua=6.51008984492044e-10 lua=-2.96739726801554e-16 wua=-2.31090391842434e-15 pua=8.64805142938968e-22 ub=-9.38661973593503e-19 lub=1.72900451661168e-24 wub=2.15724513182886e-24 pub=-1.36673579945642e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0339759495312918 lu0=6.68201910543191e-09 wu0=-3.70066788952102e-09 pu0=-4.05072860921851e-15 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.909235054012761+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.5081503516459e-08 wnfactor=3.50597320194698e-08 pnfactor=2.87812885803869e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.71063153745687 lpclm=1.11202699939703e-06 wpclm=8.72349941272644e-06 ppclm=-3.23852064547998e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.55004225855407e-05 lalpha0=-4.09605883407871e-12 walpha0=1.94829314550073e-11 palpha0=-7.23286295628836e-18 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960162e-8 kt2=-0.019151 at=-3178.99199999991 lat=0.019593725769072 ute=-1.300956205 lute=8.74719900405075e-10 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=7.97979572520804e-18 lub1=-4.28126099732196e-24 wub1=-5.5954439818879e-24 pub1=2.07725821928005e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.48 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.78279975596+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=2.89137074138829e-8 k1=0.88325 k2=-0.041769513184 wk2=8.03935420934133e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=42099.668128 wvsat=0.104621282132206 ua=-1.473525560832e-10 wua=2.66954817810876e-18 ub=1.64936923264e-18 wub=3.76412873757972e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.040807699868 wu0=-2.88314493558059e-9 a0=0.8137278731976 wa0=4.27228337521772e-7 keta=-0.034899157736 wketa=1.33066118615052e-8 a1=0.0 a2=0.65972622 ags=0.1523008606664 wags=5.06992057083846e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.05908438768+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=-1.31996763860058e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.33242727464 wpclm=-1.26120796578128e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=21.0696152 wbeta0=7.95161228072641e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414028144 wkt1=3.29032232305917e-8 kt2=-0.019151 at=154649.9232 wat=-0.119548377737818 ute=-1.407344636 wute=3.16693523594449e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.49 nmos lmin=8e-06 lmax=2.0e-05 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.78279975596+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=2.89137074138829e-8 k1=0.88325 k2=-0.041769513184 wk2=8.0393542093413e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=42099.668128 wvsat=0.104621282132206 ua=-1.473525560832e-10 wua=2.66954817810866e-18 ub=1.64936923264e-18 wub=3.76412873757972e-25 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.040807699868 wu0=-2.88314493558061e-9 a0=0.813727873197601 wa0=4.27228337521771e-7 keta=-0.034899157736 wketa=1.33066118615052e-8 a1=0.0 a2=0.65972622 ags=0.1523008606664 wags=5.06992057083845e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.05908438768+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=-1.31996763860058e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.33242727464 wpclm=-1.26120796578128e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.4467e-5 alpha1=0.0 beta0=21.0696152 wbeta0=7.95161228072641e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.414028144 wkt1=3.29032232305919e-8 kt2=-0.019151 at=154649.9232 wat=-0.119548377737818 ute=-1.407344636 wute=3.16693523594448e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.50 nmos lmin=4e-06 lmax=8e-06 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.775077003430057+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=6.07876463465396e-08 wvth0=3.98203036838399e-08 pvth0=-8.58484477305355e-14 k1=0.88325 k2=-0.0443174578143169 lk2=2.00554862398803e-08 wk2=1.16377348765097e-08 pk2=-2.83237214410232e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=27007.4179283649 lvsat=0.118794738553626 wvsat=0.125935584137144 pvsat=-1.67770007827653e-7 ua=-1.483548227984e-10 lua=7.88908286161658e-18 wua=4.08501738745059e-18 pua=-1.11414992748094e-23 ub=1.36246239959938e-18 lub=2.25831282740951e-24 wub=7.81602213042588e-25 pub=-3.18934294013998e-30 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0397702955682965 lu0=8.16565925740254e-09 wu0=-1.41805204004695e-09 pu0=-1.15320992681334e-14 a0=0.822752031664827 la0=-7.10313261177352e-08 wa0=4.14483807291578e-07 pa0=1.00315268873639e-13 keta=-0.034899157736 wketa=1.33066118615052e-8 a1=0.0 a2=0.65972622 ags=0.103616891779771 lags=3.83203251943161e-07 wags=1.19454017079967e-07 pags=-5.41185690215264e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.18169013039989+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-9.65059348932287e-07 wnfactor=-3.05148930919598e-07 pnfactor=1.3629224365979e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.33242727464 wpclm=-1.26120796578128e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.55549498089627e-05 lalpha0=-8.56351514224969e-12 walpha0=-1.5364767008042e-12 palpha0=1.20939784029147e-17 alpha1=0.0 beta0=15.6204710791158 lbeta0=4.28915266192126e-05 wbeta0=1.56472641500393e-05 pbeta0=-6.05743305154622e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.436576326569176 lkt1=1.77482179113983e-07 wkt1=6.47472999311968e-08 pkt1=-2.50652402132948e-13 kt2=-0.019151 at=255365.138675653 lat=-0.792753733375793 wat=-0.261785253667187 pat=1.11958072952716e-6 ute=-1.48250524456392 lute=5.91607263713278e-07 wute=4.22840445929798e-07 pute=-8.35508007109826e-13 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.51 nmos lmin=2e-06 lmax=4e-06 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.787310399081536+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.34292235313137e-08 wvth0=1.69132113658525e-08 pvth0=2.83042724164143e-15 k1=0.88325 k2=-0.0439173137240638 lk2=1.85064320317849e-08 wk2=5.83744779518737e-09 pk2=-5.86941228003773e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=27734.1731690256 lvsat=0.115981293869016 wvsat=0.131582012773011 pvsat=-1.89628693866396e-7 ua=-1.45545872992138e-10 lua=-2.98503879532675e-18 wua=3.38862529026679e-18 pua=-8.4455976361154e-24 ub=1.99792193506897e-18 lub=-2.01704180141344e-25 wub=-9.32022819309903e-26 pub=1.97236087786037e-31 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0409046390641042 lu0=3.77434220834841e-09 wu0=-4.48542276373835e-09 pu0=3.4243203962045e-16 a0=0.514935664325726 la0=1.12060001559645e-06 wa0=8.54915327510911e-07 pa0=-1.60470128989177e-12 keta=-0.0272934850239557 lketa=-2.94433920354469e-08 wketa=-8.84314539625447e-09 pketa=8.5747048436287e-14 a1=0.0 a2=0.65972622 ags=0.20819955184146 lags=-2.16614295767118e-08 wags=-3.67251314347774e-08 pags=6.34214328601026e-14 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.953883122762372+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-8.31635208785952e-08 wnfactor=2.89566365234256e-08 pnfactor=6.95192655842022e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.33242727464 wpclm=-1.26120796578128e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.12719014791517e-05 lalpha0=8.01719715709617e-12 walpha0=6.04113375222549e-12 palpha0=-1.72407778648824e-17 alpha1=0.0 beta0=22.7625727189021 lbeta0=1.52427299251048e-05 wbeta0=2.74755501772768e-06 pbeta0=-1.06364476343831e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207288e-8 kt2=-0.019151 at=97365.905 lat=-0.181100622002025 wat=0.02741935269216 ute=-1.26724183483923 lute=-2.41729273812727e-07 wute=1.34158444755344e-07 pute=2.82049591798768e-13 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.52 nmos lmin=1e-06 lmax=2e-06 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.782033376158791+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=2.33038051822929e-08 wvth0=1.45796978634537e-08 pvth0=7.19699338138591e-15 k1=0.88325 k2=-0.0402352415445912 lk2=1.16163876045962e-08 wk2=6.38241700066917e-10 pk2=3.85955533260156e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=81477.7326095998 lvsat=0.015414141957876 wvsat=0.0516957461239179 pvsat=-4.01422363756798e-8 ua=-1.48488361317388e-10 lua=2.52106600090287e-18 wua=-7.23647816526074e-19 pua=-7.50543595487271e-25 ub=1.83194351969081e-18 lub=1.08881435829302e-25 wub=1.31137100433649e-25 pub=-2.22556962409352e-31 uc=6.6204e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0422333031731971 lu0=1.28809145218538e-09 wu0=-4.11184011057494e-09 pu0=-3.56631137867635e-16 a0=1.13092924284003 la0=-3.20724242562321e-08 wa0=-1.57273330785289e-08 pa0=2.44809529522735e-14 keta=-0.0712286511851589 lketa=5.2769892227209e-08 wketa=6.91993922018543e-08 pketa=-6.02893476613358e-14 a1=0.0 a2=0.65972622 ags=0.151565191558124 lags=8.43151073942377e-08 wags=3.61948184066163e-08 pags=-7.3029367001056e-14 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.948201532380995+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.25318960117566e-08 wnfactor=4.20041953035985e-08 pnfactor=4.5104138644834e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.92049697412599 lpclm=-1.10042013253586e-06 wpclm=-2.97382453336394e-06 ppclm=3.20471833853995e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.00821580576818e-05 lalpha0=-8.46891617316897e-12 walpha0=-2.73646719414407e-11 palpha0=4.52695353871393e-17 alpha1=0.0 beta0=29.4253813627996 lbeta0=2.77500921548936e-06 wbeta0=-9.02827305934221e-06 pbeta0=1.13989646723812e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=-19815.33256392 lat=0.0381737141583222 wat=0.0513082169510301 pat=-4.47018222446325e-8 ute=-1.48165058947913 lute=1.59481178628385e-07 wute=5.33092374121203e-07 pute=-4.64451933121731e-13 ua1=3.0044e-9 ub1=-4.2599574569176e-18 lub1=9.49575199139945e-25 wub1=7.16665927766103e-25 pub1=-1.34105466733897e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.53 nmos lmin=8.0e-07 lmax=1e-06 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.824404809240084+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.36119245468858e-08 wvth0=-6.58616261933963e-08 pvth0=7.72807729940001e-14 k1=0.88325 k2=-0.0240682856376772 lk2=-2.46892722669942e-09 wk2=-1.77070663277373e-08 pk2=1.98427398440538e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=97530.4993496758 lvsat=0.00142831341048544 wvsat=-0.0518661103342097 pvsat=5.00850990067556e-8 ua=-1.32089692140148e-10 lua=-1.17661269317445e-17 wua=-6.69762149684785e-17 pua=5.6971409262547e-23 ub=1.18219860440148e-19 lub=1.60194775043851e-24 wub=2.06462239136185e-24 pub=-1.90708862076293e-30 uc=6.4949516809062e-11 luc=1.09295718975609e-18 wuc=3.65339125350693e-18 puc=-3.18298424909669e-24 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0337284867791748 lu0=8.69783619212973e-09 wu0=1.53206945147825e-08 pu0=-1.72870520373987e-14 a0=0.999864250024796 la0=8.21167711491053e-08 wa0=5.38932777680129e-08 pa0=-3.61753776622781e-14 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.543992731012645 lags=-2.57583854507659e-07 wags=-2.07474786088287e-07 pags=1.39265582888688e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.08601980340374+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.92604824275881e-07 wnfactor=-4.08314042486365e-07 pnfactor=4.37439850455201e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.720234099675163 lpclm=-5.47019055364481e-08 wpclm=1.22491404551775e-06 ppclm=-4.53394859663518e-13 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.55853129544524e-05 lalpha0=-4.55108034858631e-12 walpha0=-4.7608056192314e-12 palpha0=2.55761202887113e-17 alpha1=0.0 beta0=27.643516649718 lbeta0=4.32744280997921e-06 wbeta0=4.06452476003064e-06 pbeta0=-8.01759256693041e-15 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37944241 lkt1=5.84812680081025e-9 kt2=-0.019151 at=7218.97500000001 lat=0.014620317002025 ute=-1.4714445575 lute=1.50589265120857e-7 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-1.13102438357546e-17 lub1=7.0920737541243e-24 wub1=1.42466915250071e-24 pub1=-1.95789610485997e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.54 nmos lmin=6e-07 lmax=8.0e-07 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.728980208989632+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=5.04409795498282e-08 wvth0=7.43494607552888e-08 pvth0=-1.68346572205225e-14 k1=0.88325 k2=-0.0214639589703167 lk2=-4.21705806322515e-09 wk2=-1.67097694136341e-09 pk2=9.07865916825475e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=89724.2801147174 lvsat=0.00666816781597807 wvsat=0.0528454428506869 pvsat=-2.02015886646277e-8 ua=-1.50831218484322e-10 lua=8.13953953044598e-19 wua=1.16414769559746e-17 pua=4.19999111748507e-24 ub=2.81006265736214e-18 lub=-2.04927500410208e-25 wub=-3.29264638547404e-24 pub=1.68892983026917e-30 uc=5.21848316746435e-11 luc=9.66113720406823e-18 wuc=4.08275753005493e-17 puc=-2.81358207230174e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0497666263024752 lu0=-2.06762061962997e-09 wu0=-2.50951207217259e-08 pu0=9.84170019777039e-15 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.723635362438653+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=5.06424702619624e-08 wnfactor=7.10601988756954e-07 pnfactor=-3.13622465272598e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.142499392724535 lpclm=3.33097316891797e-07 wpclm=-1.14392139001962e-06 ppclm=1.13666460692202e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-1.01867832456375e-05 lalpha0=1.27482072768582e-11 walpha0=1.02553929198083e-10 palpha0=-4.64579296247974e-17 alpha1=0.0 beta0=27.3291860472631 lbeta0=4.53843439790169e-06 wbeta0=1.36012903594039e-05 pbeta0=-6.40948567025583e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67299999998 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210592e-8 ua1=2.0117e-9 ub1=4.26468502581761e-19 lub1=-7.86088772572957e-25 wub1=-3.14606494080414e-24 pub1=1.11016801866406e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.55 nmos lmin=5e-07 lmax=6e-07 wmin=1.5e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.802305943849357+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.58868869287956e-08 wvth0=-3.02989313323749e-08 pvth0=3.24799557152605e-14 k1=0.88325 k2=-0.0242385648208956 lk2=-2.9095500275925e-09 wk2=6.59011097700796e-08 pk2=-2.27640785457324e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=86072.415023637 lvsat=0.00838907637336389 wvsat=-0.00968864165167704 pvsat=9.2670358503509e-9 ua=-1.69630873270131e-10 lua=9.67312207396408e-18 wua=7.90192788609986e-17 pua=-2.75511916300403e-23 ub=-1.86461676764022e-18 lub=1.99797310650733e-24 wub=4.85387364797769e-24 pub=-2.15004441681466e-30 uc=9.67513030325892e-11 luc=-1.13404113251214e-17 wuc=-8.89619331081125e-17 puc=3.30263170089888e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.031115656533084 lu0=6.72148102546771e-09 wu0=4.62927187978349e-09 pu0=-4.16565229615741e-15 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.16818579371347+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.58847919522416e-07 wnfactor=-7.19074220787247e-07 pnfactor=3.60099581389222e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.767215635813001 lpclm=7.61792336654854e-07 wpclm=5.97601947167785e-06 ppclm=-2.21854344468516e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.57703380640077e-05 lalpha0=-4.1962625262203e-12 walpha0=1.86968652443629e-11 palpha0=-6.94104295018255e-18 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960162e-8 kt2=-0.019151 at=-3178.99200000003 lat=0.019593725769072 ute=-1.300956205 lute=8.74719900405075e-10 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=6.63808752273775e-18 lub1=-3.71325833125028e-24 wub1=-1.68803011849615e-24 pub1=4.23082230964826e-31 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.56 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.799704207584+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=5.04009132775877e-9 k1=0.88325 k2=-0.036365276688 wk2=4.07123941608392e-10 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123989.01408 wvsat=-0.0110284206967335 ua=-1.464891488608e-10 wua=1.45018578694419e-18 ub=2.15693945096e-18 wub=-3.40412303328377e-25 uc=9.0941059088e-11 wuc=-3.49353569640916e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0416743279304 wu0=-4.10705601601016e-9 a0=1.1105683473904 wa0=8.01003471445444e-9 keta=-0.032116486504 wketa=9.37673432603107e-9 a1=0.0 a2=0.65972622 ags=0.218854029336 wags=-4.32917047022941e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.804476980479999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=2.27577129891471e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.634185227760002 wpclm=1.51617593975816e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-1.5360514528e-05 walpha0=4.21244442874296e-11 alpha1=0.0 beta0=26.214673424 wbeta0=6.85411192834391e-7 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.387080928 wkt1=-5.15346761529579e-9 kt2=-0.019151 at=-75962.8800000003 wat=0.20613870461184 ute=-1.2093733184 wute=3.71049668301313e-8 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.57 nmos lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.799704207584+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=5.04009132775962e-9 k1=0.88325 k2=-0.036365276688 wk2=4.07123941608392e-10 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123989.01408 wvsat=-0.0110284206967334 ua=-1.464891488608e-10 wua=1.45018578694429e-18 ub=2.15693945096e-18 wub=-3.4041230332838e-25 uc=9.0941059088e-11 wuc=-3.49353569640916e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0416743279304 wu0=-4.10705601601018e-9 a0=1.1105683473904 wa0=8.01003471445487e-9 keta=-0.032116486504 wketa=9.37673432603107e-9 a1=0.0 a2=0.65972622 ags=0.218854029336 wags=-4.32917047022942e-8 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.804476980479999+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=2.27577129891471e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.634185227760001 wpclm=1.51617593975816e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-1.5360514528e-05 walpha0=4.21244442874296e-11 alpha1=0.0 beta0=26.214673424 wbeta0=6.85411192834378e-7 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.387080928 wkt1=-5.15346761529579e-9 kt2=-0.019151 at=-75962.8800000002 wat=0.20613870461184 ute=-1.2093733184 wute=3.71049668301309e-8 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.58 nmos lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.810194852963869+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-8.25743980304825e-08 wvth0=-9.77551144157701e-09 pvth0=1.16617179957712e-13 k1=0.88325 k2=-0.0327697452753609 lk2=-2.83012942719525e-08 wk2=-4.67073001545653e-09 pk2=3.99690122588616e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123989.01408 wvsat=-0.0110284206967335 ua=-1.4005455674428e-10 lua=-5.06482252858237e-17 wua=-7.63718275226833e-18 pua=7.15288678279601e-23 ub=3.00752754715302e-18 lub=-6.69518389686644e-24 wub=-1.5416706527627e-24 pub=9.45539397165978e-30 uc=9.0941059088e-11 wuc=-3.49353569640916e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0439348580593255 lu0=-1.77931774325339e-08 wu0=-7.29953038012751e-09 pu0=2.51287351062897e-14 a0=1.09536176755236 la0=1.19694654690977e-07 wa0=2.94858008091685e-08 pa0=-1.6904093059112e-13 keta=-0.032116486504 wketa=9.37673432603109e-9 a1=0.0 a2=0.65972622 ags=0.306344351947741 lags=-6.88657414444762e-07 wags=-1.66851487636532e-07 pags=9.72568829383076e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.744580887013387+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.71456586634237e-07 wnfactor=3.12166466019378e-07 pnfactor=-6.65823050692758e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.634185227760001 wpclm=1.51617593975816e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-3.14540580378675e-05 lalpha0=1.26676159510153e-10 walpha0=6.48528407930231e-11 palpha0=-1.78900686439085e-16 alpha1=0.0 beta0=28.1994378419384 lbeta0=-1.56225590618183e-05 wbeta0=-2.11760808215873e-06 pbeta0=2.2063240241116e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.383549318715412 lkt1=-2.77981477968303e-08 wkt1=-1.01410463964226e-08 pkt1=3.92584345927327e-14 kt2=-0.019151 at=-270201.39065234 lat=1.52889812882564 wat=0.480455537573799 pat=-2.15921390260032e-6 ute=-1.2093733184 wute=3.71049668301317e-8 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.59 nmos lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.7709994544538+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=6.91604356930346e-08 wvth0=3.99486365133757e-08 pvth0=-7.58769802955668e-14 k1=0.88325 k2=-0.0416469968279836 lk2=6.06468590587393e-09 wk2=2.63115189299387e-09 pk2=1.17016676377101e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=134091.178451452 lvsat=-0.0391079129035048 wvsat=-0.0186225823631909 pvsat=2.93988300038181e-8 ua=-1.48483561197971e-10 lua=-1.80175176555144e-17 wua=7.53742833734271e-18 pua=1.27842912188034e-23 ub=5.83006262229867e-19 lub=2.69072230670075e-24 wub=1.90503784551815e-24 pub=-3.88764528193347e-30 uc=1.13407850586463e-10 luc=-8.69743643873003e-17 wuc=-6.66644876600426e-17 puc=1.22831111644524e-22 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0368299040003206 lu0=9.71181202380253e-09 wu0=1.26919517532121e-09 pu0=-8.04286658171124e-15 a0=1.14188715098701 la0=-6.04163172019607e-08 wa0=-3.05081946532426e-08 pa0=6.32102843967785e-14 keta=-0.0549335046401328 lketa=8.83301761063409e-08 wketa=3.01919698270447e-08 pketa=-8.05807930961795e-14 a1=0.0 a2=0.65972622 ags=0.0569997420438959 lags=2.76615662544009e-07 wags=1.76809521548408e-07 pags=-3.57825759475043e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.764479515378006+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.94424200665359e-07 wnfactor=2.96445290316929e-07 pnfactor=-6.04962590745234e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.634185227760001 wpclm=1.51617593975816e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-7.03466942416486e-06 lalpha0=3.21428211138541e-11 walpha0=3.18949180287106e-11 palpha0=-5.1312624559045e-17 alpha1=0.0 beta0=21.0606542072332 lbeta0=1.20133928349816e-05 wbeta0=5.15112007036525e-06 pbeta0=-6.07575820078903e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=222729.30353764 lat=-0.379355384681077 wat=-0.149627363433796 pat=2.7998885717922e-7 ute=-1.17871807049878 lute=-1.1867385254037e-07 wute=9.13916513778106e-09 pute=1.08262358109299e-13 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.60 nmos lmin=1e-06 lmax=2e-06 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.802094037382234+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.09749772394509e-08 wvth0=-1.37513320412537e-08 pvth0=2.46086025625674e-14 k1=0.88325 k2=-0.0516094978765278 lk2=2.47069263304528e-08 wk2=1.67017399414583e-08 pk2=-1.46277936126866e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=129014.255836002 lvsat=-0.0296077671516475 wvsat=-0.0154385644599868 pvsat=2.34407651586086e-8 ua=-1.70643556464263e-10 lua=2.34491740465779e-17 wua=3.05654253231612e-17 pua=-3.03066408889366e-23 ub=2.04807649563215e-18 lub=-5.07771819211676e-26 wub=-1.7410058523307e-25 pub=2.9237943638685e-33 uc=3.59881606735583e-11 luc=5.7896533585013e-17 wuc=4.26728629738752e-17 puc=-8.17654216930391e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0424824498995604 lu0=-8.65463617236893e-10 wu0=-4.46370205952266e-09 pu0=2.6847657729152e-15 a0=1.10298758182593 la0=1.23741514945792e-08 wa0=2.37337806385311e-08 pa0=-3.82895236901744e-14 keta=-0.00517622098996585 lketa=-4.77769310848115e-09 wketa=-2.40843412850505e-08 pketa=2.09832655855287e-14 a1=0.0 a2=0.65972622 ags=0.218087937662943 lags=-2.48191737143721e-08 wags=-5.77531271893444e-08 pags=8.10974859116379e-14 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.08384367973116+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.03183117603003e-07 wnfactor=-1.49558868850326e-07 pnfactor=2.29618678059059e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-2.39839432621797 lpclm=3.30126039760759e-06 wpclm=3.12560744559022e-06 ppclm=-3.01163422040468e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-3.3820225625529e-06 lalpha0=2.53078385478845e-11 walpha0=5.77303949473688e-12 palpha0=-2.43229444925346e-18 alpha1=0.0 beta0=20.5095793123789 lbeta0=1.30445867723037e-05 wbeta0=3.56322887080126e-06 pbeta0=-3.10443108462577e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=16515.036 lat=0.00652120752032402 ute=-0.862624794623803 lute=-7.10160550181936e-07 wute=-3.41137947127538e-07 pute=7.63715251941764e-13 ua1=3.0044e-9 ub1=-3.03669836070005e-18 lub1=-1.33943737532529e-24 wub1=-1.01090374953087e-24 pub1=1.89164454317589e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.61 nmos lmin=8.0e-07 lmax=1e-06 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.733061652267425+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=7.1118821479261e-08 wvth0=6.31393914180681e-08 pvth0=-4.23817482348554e-14 k1=0.88325 k2=-0.0363352925414555 lk2=1.13994124001192e-08 wk2=-3.82765021752156e-10 pk2=2.56927575965946e-16 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=25436.261971334 lvsat=0.0606336278009998 wvsat=0.0499502740996265 pvsat=-3.35286719369074e-8 ua=-1.66496949929517e-10 lua=1.98364804226393e-17 wua=-1.83839458248018e-17 pua=1.23400581793858e-23 ub=2.10680932039939e-18 lub=-1.01947626904209e-25 wub=-7.43798868075876e-25 pub=4.99268296006118e-31 uc=2.25392690957023e-10 luc=-1.07120458783683e-16 wuc=-2.22935369414086e-16 puc=1.4964336030088e-22 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0488401135245301 lu0=-6.40452083151905e-09 wu0=-6.02097236562688e-09 pu0=4.04152351167572e-15 a0=1.10037752536093 la0=1.46481396992054e-08 wa0=-8.80584045643979e-08 pa0=5.91084115382115e-14 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.288108044665139 lags=-8.58235617590727e-08 wags=1.53902968130332e-07 pags=-1.03305982230772e-13 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.445278569798267+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.53160987340041e-07 wnfactor=4.96584298015162e-07 pnfactor=-3.33327740783995e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=2.60889713319558 lpclm=-1.06129722078334e-06 wpclm=-1.44238431950607e-06 ppclm=9.68187493009572e-13 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=3.01838027231681e-06 lalpha0=1.97315451816298e-11 walpha0=1.29870712659029e-11 palpha0=-8.71745470359595e-18 alpha1=0.0 beta0=30.52152901 lbeta0=4.32176570579863e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37944241 lkt1=5.84812680081025e-9 kt2=-0.019151 at=7218.97500000003 lat=0.014620317002025 ute=-3.12304993887387 lute=1.25921451291963e-06 wute=2.33250942874211e-06 pute=-1.56567596145828e-12 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-1.38804710129998e-17 lub1=8.10810195403697e-24 wub1=5.05451874765433e-24 pub1=-3.39280021869424e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.62 nmos lmin=6e-07 lmax=8.0e-07 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.781625642260999+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.85206802719842e-8 k1=0.88325 k2=-0.022647145831 lk2=2.21136711404626e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=127143.128981 lvsat=-0.00763619131743531 ua=-1.42588110975e-10 lua=3.78788745397006e-18 ub=4.78602633149995e-19 lub=9.90971458051762e-25 uc=8.10940580400001e-11 luc=-1.02613001258276e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0319972505737 lu0=4.90109933845903e-9 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.22679905995+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.71427607989898e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.6674894975 lpclm=1.1379478175914e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=6.2429695495e-05 lalpha0=-2.01477654597593e-11 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67300000001 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210592e-8 ua1=2.0117e-9 ub1=-1.8012e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.63 nmos lmin=5e-07 lmax=6e-07 wmin=1e-06 wmax=1.5e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.753521076540748+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=5.17647039265613e-08 wvth0=3.8598375651822e-08 pvth0=-1.81891371405406e-14 k1=0.88325 k2=0.0415632699551387 lk2=-2.80472134314295e-08 wk2=-2.70287158254008e-08 pk2=1.27370390742777e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=92324.7476956779 lvsat=0.00877165749784081 wvsat=-0.018518611009755 pvsat=8.72672877084804e-9 ua=-4.96699581928675e-11 lua=-3.99989557812348e-17 wua=-9.03976827533374e-17 pua=4.25990944183656e-23 ub=1.03017347323152e-18 lub=7.31048663800903e-25 wub=7.65654024082235e-25 pub=-3.60807567962537e-31 uc=-1.00767950514046e-10 luc=7.54395346471894e-17 wuc=1.89988188059686e-16 puc=-8.95302237294348e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0285257368668284 lu0=6.53701892919897e-09 wu0=8.28693254700701e-09 pu0=-3.90514238038414e-15 a0=1.1222 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.705217833717803+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.43628506409882e-08 wnfactor=-6.52393858600813e-08 pnfactor=3.07434734320904e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=3.464289625 lpclm=-8.09115907874626e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=3.900923128e-05 lalpha0=-9.11108248261848e-12 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.4449782 lkt1=3.49887960162e-8 kt2=-0.019151 at=-62134.8892210791 lat=0.0473761617314306 wat=0.083261527056619 pat=-3.92362452716882e-8 ute=-0.245656482223787 lute=-4.96425776760379e-07 wute=-1.49036602888571e-06 pute=7.02321577818132e-13 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=1.89429403792469e-17 lub1=-9.77548945645669e-24 wub1=-1.90657800524526e-23 pub1=8.98457725769782e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.64 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.7408250264432+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=5.87536841487147e-8 k1=0.88325 k2=-0.042411875472 wk2=5.9232425210905e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=140774.8848 wvsat=-0.0263416334067264 ua=-1.61931708424e-10 wua=1.55379387145457e-17 ub=2.58692758880001e-19 wub=1.39129740996206e-24 uc=4.1106642368e-11 wuc=1.05269867082294e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0346223032928 wu0=2.32628039608394e-9 a0=1.9441868048464 wa0=-7.52473408232016e-7 keta=-0.026034130048 wketa=3.82799516662887e-9 a1=0.0 a2=0.65972622 ags=0.200933503728 wags=-2.6943382646935e-8 b0=5.2385902304e-07 wb0=-4.47856101186655e-13 b1=-6.1646554512e-10 wb1=5.62381789915532e-16 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0747352152+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=-1.89708093800739e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=3.20594647056 wpclm=-1.98705332440483e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=3.8097298928e-05 walpha0=-6.64340827844871e-12 alpha1=0.0 beta0=22.30363328 wbeta0=4.25332796292096e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.398028144 wkt1=4.83332723059204e-9 kt2=-0.019151 at=388416.48 wat=-0.21749972537664 ute=-1.264066592 wute=8.69998901506558e-8 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.65 nmos lmin=8e-06 lmax=2.0e-05 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.698580093341266+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=8.39459246697396e-07 wvth0=9.72923847797495e-08 pvth0=-7.65811808066139e-13 k1=0.88325 k2=-0.0466707911072584 lk2=8.46299389868878e-08 wk2=9.80851496983641e-09 pk2=-7.72051851796902e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=159714.982892336 lvsat=-0.376363253756457 wvsat=-0.043620078813226 pvsat=3.43344152777896e-7 ua=-1.73103759862961e-10 lua=2.22002526607996e-16 wua=2.5729843736664e-17 pua=-2.02525800943622e-22 ub=-7.41674568894219e-19 lub=1.98785402587275e-23 wub=2.30390051133599e-24 pub=-1.81345561647488e-29 uc=3.35375536257783e-11 luc=1.50407186547076e-16 wuc=1.74320241569186e-17 puc=-1.37211663256928e-22 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0329496667401685 lu0=3.32373640427491e-08 wu0=3.85217319867996e-09 pu0=-3.03213836205506e-14 a0=2.48522843061551 la0=-1.07511685366897e-05 wa0=-1.24604837008915e-06 pa0=9.80794701862887e-12 keta=-0.0287865259542625 lketa=5.46935223807547e-08 wketa=6.33891787524311e-09 pketa=-4.98951502752464e-14 a1=0.0 a2=0.65972622 ags=0.220306270116207 lags=-3.84960909736765e-07 wags=-4.46165374943722e-08 pags=3.51187519203739e-13 b0=8.45875443083283e-07 lb0=-6.3988658886373e-12 wb0=-7.416213766667e-13 pb0=5.83748058649538e-18 b1=-1.02082795127299e-09 lb1=8.03518282400597e-15 wb1=9.31268673451909e-16 pb1=-7.33024016449028e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.08837556107384+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.71050600182408e-07 wnfactor=-3.14144604297097e-08 pnfactor=2.47270788927206e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=4.6346727874831 lpclm=-2.83905649666212e-05 wpclm=-3.29043462409163e-06 ppclm=2.58998039209696e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.28740264193608e-05 lalpha0=-9.49195031721559e-11 walpha0=-1.10010639135375e-11 palpha0=8.65920253198565e-17 alpha1=0.0 beta0=19.245415606375 lbeta0=6.07705804230607e-05 wbeta0=7.04324208360346e-06 pbeta0=-5.54390558613849e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.401503391356392 lkt1=6.90574777534787e-08 wkt1=8.00368418591313e-09 pkt1=-6.29989271152101e-14 kt2=-0.019151 at=544802.61103764 lat=-3.10758649890652 wat=-0.360165788366086 pat=2.83495172018446e-6 ute=-1.32662104441506 lute=1.24303459956262e-06 wute=1.44066315346435e-07 pute=-1.13398068807379e-12 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.66 nmos lmin=4e-06 lmax=8e-06 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.846578534989263+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-3.25472155138423e-07 wvth0=-4.29671802755193e-08 pvth0=3.38205031039057e-13 k1=0.88325 k2=-0.0368261913915029 lk2=7.14072207564472e-09 wk2=-9.70164029975967e-10 pk2=7.63639488947198e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=83954.5905229907 lvsat=0.219965052837223 wvsat=0.0254937028127722 pvsat=-2.00667078821708e-7 ua=-1.41284738340155e-10 lua=-2.84526601821995e-17 wua=-6.51492744816304e-18 pua=5.12805640420066e-23 ub=1.55861854981662e-18 lub=1.77237875071289e-24 wub=-2.19877339580618e-25 pub=1.73070753027787e-30 uc=6.38139085946653e-11 luc=-8.7905300014582e-17 wuc=-1.01881256378382e-17 puc=8.01931922337028e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0351191526928434 lu0=1.61608172631308e-08 wu0=7.42755523142404e-10 pu0=-5.84640772673486e-15 a0=0.351475087215166 la0=6.04411826377011e-06 wa0=7.08109814907017e-07 pa0=-5.57370300759852e-12 keta=-0.0177769423292126 lketa=-3.19655636416662e-08 wketa=-3.70477295921386e-09 pketa=2.91611608122555e-14 a1=0.0 a2=0.65972622 ags=-0.0321654406601031 lags=1.60230477146587e-06 wags=1.41960163846241e-07 pags=-1.11740266203325e-12 b0=-4.42190237089848e-07 lb0=3.73980950383433e-12 wb0=4.33439725253481e-13 pb0=-3.41170853644394e-18 b1=5.96621673338973e-10 lb1=-4.69615297667433e-15 wb1=-5.44278860693599e-16 pb1=4.28415008372474e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.15360636451171+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.84497974665512e-07 wnfactor=-6.09743882870609e-08 pnfactor=4.7994410503504e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.08023248020929 lpclm=1.65928316875551e-05 wpclm=1.92309057465557e-06 ppclm=-1.51371093779425e-11 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=5.59542034736526e-05 lalpha0=-1.97876729089157e-10 walpha0=-1.48869191195684e-11 palpha0=1.1717852813763e-16 alpha1=0.0 beta0=27.508757464998 lbeta0=-4.27217481154798e-06 wbeta0=-1.48752247604799e-06 pbeta0=1.17086479018904e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.3946656205 lkt1=1.52357354400412e-8 kt2=-0.019151 at=307735.10819176 lat=-1.24157105073842 wat=-0.0467774363537105 pat=3.68196474902217e-7 ute=-1.07640323475483 lute=-7.26490082765141e-07 wute=-8.41993854366791e-08 pute=6.6275365482399e-13 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.67 nmos lmin=2e-06 lmax=4e-06 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.769921428700284+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-2.87140223311684e-08 wvth0=4.09320849114852e-08 pvth0=1.34107557772552e-14 k1=0.88325 k2=-0.0439534431571026 lk2=3.47320313279568e-08 wk2=4.73524907276672e-09 pk2=-1.44506342358025e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=172047.023973194 lvsat=-0.121061987324976 wvsat=-0.0532484856456195 pvsat=1.04162909568145e-7 ua=-1.45661056358777e-10 lua=-1.15108784394717e-17 wua=4.9625474927003e-18 pua=6.84849247446335e-24 ub=2.27570496377101e-18 lub=-1.00363557553031e-24 wub=3.60842986460614e-25 pub=-5.17400805426306e-31 uc=-3.82694062892532e-12 luc=1.739487287746e-16 wuc=4.02850608524371e-17 puc=-1.15200676708097e-22 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0383435754229819 lu0=3.67829978888648e-09 wu0=-1.11678826087217e-10 pu0=-2.53868644218893e-15 a0=1.57064013617825 la0=1.32443654045721e-06 wa0=-4.21645822947687e-07 pa0=-1.20014666235424e-12 keta=-0.026034130048 wketa=3.82799516662885e-9 a1=0.0 a2=0.65972622 ags=0.490720460893236 lags=-4.2191256894938e-07 wags=-2.18860011194842e-07 pags=2.79419193212968e-13 b0=8.15871528932108e-07 lb0=-1.13045078532227e-12 wb0=-7.14249765911837e-13 pb0=1.03127407702438e-18 b1=1.95225408771331e-09 lb1=-9.94413276012927e-15 wb1=-1.78097893209005e-15 pb1=9.07171410481761e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.21084710627118+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.00609068103517e-06 wnfactor=-1.10761579092002e-07 pnfactor=6.72682319353945e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=3.20594647056 wpclm=-1.98705332440483e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.75608021378663e-05 lalpha0=-8.79590297086061e-11 walpha0=3.34576377759575e-13 palpha0=5.82524506870591e-17 alpha1=0.0 beta0=27.5504396995595 lbeta0=-4.43353678695438e-06 wbeta0=-7.69303561148297e-07 pbeta0=8.92824939155525e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=-43839.55138352 lat=0.119459185970449 wat=0.093554872707421 pat=-1.75063713559907e-7 ute=-1.35329353049034 lute=3.45418982588267e-07 wute=1.68398770873358e-07 pute=-3.15114684407832e-13 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.68 nmos lmin=1e-06 lmax=2e-06 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.698018016979329+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.05834589720965e-07 wvth0=8.1193890939663e-08 pvth0=-6.1928786396718e-14 k1=0.88325 k2=-0.0222925455606549 lk2=-5.80072835131785e-09 wk2=-1.00431775138384e-08 pk2=1.3203363508543e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=104595.148109461 lvsat=0.0051567283181525 wvsat=0.00683820610748953 pvsat=-8.27377159463484e-9 ua=-1.2601697048153e-10 lua=-4.82696973404967e-17 wua=-1.01459810181349e-17 pua=3.51201904736073e-23 ub=1.85885347001923e-18 lub=-2.23605969510733e-25 wub=-1.4784741032229e-27 pub=1.60589966760629e-31 uc=1.51012439196883e-10 luc=-1.15793067170026e-16 wuc=-6.22601055460415e-17 puc=7.66860430085587e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0389885659522823 lu0=2.471367065848e-09 wu0=-1.27634353870712e-09 pu0=-3.59318080681255e-16 a0=3.37214918920628 la0=-2.04662106144002e-06 wa0=-2.04634974060313e-06 pa0=1.84006592122325e-12 keta=-0.0394287024851496 lketa=2.50644731218642e-08 wketa=7.16310150359775e-09 pketa=-6.24078771709602e-15 a1=0.0 a2=0.65972622 ags=0.140292290106213 lags=2.338229917823e-07 wags=1.32173526159384e-08 pags=-1.54853485121681e-13 b0=2.92451618155391e-08 lb0=3.41516724507304e-13 wb0=3.36429676486182e-15 pb0=-3.11554779232829e-19 b1=-5.58179873186972e-09 lb1=4.1538957720401e-15 wb1=5.09209636552532e-15 pb1=-3.78946618816748e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.495094247078454+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.33255414953481e-07 wnfactor=3.87538398576895e-07 pnfactor=-2.59757029159179e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=5.69678787527362 lpclm=-4.66096456099773e-06 wpclm=-4.25936823100012e-06 ppclm=4.25204881813228e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-6.35979406094325e-05 lalpha0=8.26209472285921e-11 walpha0=6.07060946195277e-11 palpha0=-5.47172094791853e-17 alpha1=0.0 beta0=16.2066023848891 lbeta0=1.67935166935869e-05 wbeta0=7.48869702648855e-06 pbeta0=-6.52445988605492e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=16515.036 lat=0.00652120752032399 ute=-1.71616794664955 lute=1.02444446795644e-06 wute=4.37522157084682e-07 pute=-8.18709398745298e-13 ua1=3.0044e-9 ub1=-4.49170923709431e-18 lub1=1.38323863202959e-24 wub1=3.16456112655571e-25 pub1=-5.92165652701722e-31 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.69 nmos lmin=8.0e-07 lmax=1e-06 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.781013131604446+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.35258430598603e-08 wvth0=1.93947912662365e-08 pvth0=-8.08687699814447e-15 k1=0.88325 k2=-0.0528446523631309 lk2=2.08175197313782e-08 wk2=1.4678195644048e-08 pk2=-8.33491036290708e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=111335.236930446 lvsat=-0.000715513406331025 wvsat=-0.0284126119883723 pvsat=2.2438186414022e-8 ua=-3.05901119481352e-10 lua=1.08452748518257e-16 wua=1.08790017123911e-16 pua=-6.85017274836671e-23 ub=7.65469044287747e-19 lub=7.28995370947985e-25 wub=4.79862942931944e-25 pub=-2.58774410758505e-31 uc=-1.93241603001466e-10 luc=1.84135168808906e-16 wuc=1.58971300666837e-16 puc=-1.16059828571756e-22 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0464464616500472 lu0=-4.02625743976843e-09 wu0=-3.83732035739621e-09 pu0=1.87190992381017e-15 a0=0.690334600566267 la0=2.898857625813e-07 wa0=2.86010634352182e-07 pa0=-1.91982064213194e-13 keta=0.0443102156354136 lketa=-4.78923056404134e-08 wketa=-5.01475686772875e-08 pketa=4.36906178819687e-14 a1=0.0 a2=0.65972622 ags=1.24242508328364 lags=-7.26400285078391e-07 wags=-7.16689928056087e-07 pags=4.81071663998296e-13 b0=1.72445164339818e-06 lb0=-1.13541666571324e-12 wb0=-1.54311832977557e-12 pb0=1.03580429079688e-18 b1=-3.54598068456401e-09 lb1=2.38020762068743e-15 wb1=3.23488470714584e-15 pb1=-2.17138724570928e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.625349444301788+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.19771746669426e-07 wnfactor=3.32311401473585e-07 pnfactor=-2.11641004975894e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.25247158564762 lpclm=1.39351520099475e-06 wpclm=2.08021879889558e-06 ppclm=-1.27125932538108e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.622192261482e-05 lalpha0=4.36619977323116e-12 walpha0=-8.18077789980779e-12 palpha0=5.2998582214331e-18 alpha1=0.0 beta0=30.52152901 lbeta0=4.32176570579857e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37944241 lkt1=5.84812680080982e-9 kt2=-0.019151 at=7218.97500000003 lat=0.014620317002025 ute=1.83176620524772 lute=-2.06666123047669e-06 wute=-2.18761078542341e-06 pute=1.46841405121839e-12 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-6.60541663102848e-18 lub1=3.22478717562819e-24 wub1=-1.58228056327785e-24 pub1=1.06209158757519e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.70 nmos lmin=6e-07 lmax=8.0e-07 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.777954270939883+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.55790757512027e-08 wvth0=3.34927457237261e-09 pvth0=2.6835316729635e-15 k1=0.88325 k2=-0.0214579613621218 lk2=-2.50514122830131e-10 wk2=-1.08485493705456e-09 pk2=2.24589547220275e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=173909.611166514 lvsat=-0.0427179989429239 wvsat=-0.0426635651704147 pvsat=3.20040104788892e-8 ua=-1.59092930237662e-10 lua=9.90907276213283e-18 wua=1.50568184591098e-17 pua=-5.58416147870707e-24 ub=-1.40259427867709e-18 lub=2.18428836391822e-24 wub=1.71615574435867e-24 pub=-1.08862482708099e-30 uc=1.66841632926662e-10 luc=-5.75674625587264e-17 wuc=-7.82247686467057e-17 puc=4.31558981903358e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0298706344972628 lu0=7.10011735409371e-09 wu0=1.94004379481911e-09 pu0=-2.00609376708703e-15 a0=1.1222 keta=-0.0270386823616 wketa=1.49417478006521e-8 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.66716838018203+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.79539837669765e-07 wnfactor=-4.01734839029436e-07 pnfactor=2.81080927545592e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-5.36267688842133 lpclm=4.15245351863388e-06 wpclm=4.28326921074102e-06 ppclm=-2.75003708687863e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=6.1625011543175e-05 lalpha0=-1.93978050421268e-11 walpha0=7.34087419363556e-13 palpha0=-6.84164890272808e-19 alpha1=0.0 beta0=34.7129675909665 lbeta0=1.50830028127212e-06 wbeta0=2.0498957617243e-06 pbeta0=-1.37597408099558e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67300000001 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210601e-8 ua1=2.0117e-9 ub1=-1.8012e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.71 nmos lmin=5e-07 lmax=6e-07 wmin=7.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.698211302820752+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=7.31572317906307e-08 wvth0=8.90557123038129e-08 pvth0=-3.77048557500391e-14 k1=0.88325 k2=0.0325590384876379 lk2=-2.57055391490307e-08 wk2=-1.88144435930068e-08 pk2=1.06008045600224e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-3467.94588173623 lvsat=0.0408695784180504 wvsat=0.0688699979747254 pvsat=-2.05551773511897e-8 ua=-9.69085190347822e-11 lua=-1.93947713575232e-17 wua=-4.73034553312058e-17 pua=2.38025563025151e-23 ub=7.24580107411366e-18 lub=-1.89119011052625e-24 wub=-4.90466413611932e-24 pub=2.03137695421534e-30 uc=-4.35315728186549e-11 luc=4.15690172899026e-17 wuc=1.37773272252268e-16 puc=-5.86312346009374e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0338982762762993 lu0=5.20212741449881e-09 wu0=3.38573676500773e-09 pu0=-2.68736356805166e-15 a0=1.1222 keta=-0.0878430665476272 lketa=2.86535188082077e-08 wketa=7.04116417532709e-08 pketa=-2.6139688296126e-14 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.293967985175604+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.67568489673459e-07 wnfactor=3.09930690969814e-07 pnfactor=-5.42850484767842e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=11.4836986225732 lpclm=-3.78624932354271e-06 wpclm=-7.31585020739814e-06 ppclm=2.71594354684469e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.27168347549054e-05 lalpha0=-1.04874969042459e-11 walpha0=-3.38232800684504e-12 palpha0=1.25565883158915e-18 alpha1=0.0 beta0=41.4540648180672 lbeta0=-1.66838111712408e-06 wbeta0=-4.09979152344849e-06 pbeta0=1.52201070495656e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.444978199999999 lkt1=3.49887960162e-8 kt2=-0.019151 at=29133.8246399999 lat=0.00436660174282177 ute=-1.87934968299999 lute=2.73437440866603e-7 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=-4.31566122590644e-18 lub1=1.18491722255738e-24 wub1=2.15229791667743e-24 pub1=-1.01425102255299e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.72 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.8295409+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' k1=0.88325 k2=-0.033468 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=101000.0 ua=-1.3847e-10 ub=2.3595e-18 uc=5.7002e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0381349 a0=0.80798 keta=-0.020254 a1=0.0 a2=0.65972622 ags=0.16025 b0=-1.52387e-7 b1=2.3271e-10 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.04609+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.20557 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.8066e-5 alpha1=0.0 beta0=28.726 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.39073 kt2=-0.019151 at=60000.0 ute=-1.1327 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.73 nmos lmin=8e-06 lmax=2.0e-05 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.845487968672323+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-3.16888044831317e-7 k1=0.88325 k2=-0.0318602990257499 lk2=-3.1947013515255e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=93850.2894249996 lvsat=0.142073621916072 ua=-1.34252654665875e-10 lua=-8.38038855146217e-17 ub=2.7371293463425e-18 lub=-7.50396374984434e-24 uc=5.98592604829999e-11 luc=-5.67773116574676e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.03876630471555 lu0=-1.254679527123e-8 a0=0.603741826870273 la0=4.05846595966049e-6 keta=-0.0192149961879999 lketa=-2.06462951481708e-8 a1=0.0 a2=0.65972622 ags=0.152936961174249 lags=1.45319156948838e-7 b0=-2.7394519851e-07 lb0=2.41551225811805e-12 b1=3.853530410925e-10 lb1=-3.03320665652197e-15 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0409408965125+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.02319076334046e-07 wnfactor=-1.6940658945086e-21 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.333760873952502 lpclm=1.07171737750507e-05 ppclm=-3.23117426778526e-27 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.62628298742499e-05 lalpha0=3.58312281327777e-11 alpha1=0.0 beta0=29.8804486799999 lbeta0=-2.2940327942411e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.389418126500001 lkt1=-2.60685544800073e-8 kt2=-0.019151 at=965.692499999888 lat=1.17308495160061 ute=-1.109086277 lute=-4.69233980640241e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.74 nmos lmin=4e-06 lmax=8e-06 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.781699693983022+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.85204838222365e-7 k1=0.88325 k2=-0.03829110292275 lk2=1.86713937817693e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=122449.131725 lvsat=-0.0830347581482211 ua=-1.51122036002375e-10 lua=4.89790805058725e-17 ub=1.2266119609725e-18 lub=4.38568262509288e-24 uc=4.8430218551e-11 luc=3.31834317884081e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0362406858533499 lu0=7.33295946729128e-9 a0=1.42069451938918 la0=-2.37196556875465e-6 keta=-0.023371011436 lketa=1.20667024685121e-8 a1=0.0 a2=0.65972622 ags=0.18218911647725 lags=-8.49316072105078e-8 b0=2.1228759553e-07 lb0=-1.41174324587415e-12 pb0=-3.85185988877447e-34 b1=-2.252191232775e-10 lb1=1.77275399712591e-15 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.0615373104625+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.9800261602164e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.8235626218575 lpclm=-6.26363937543226e-6 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=3.34755103772501e-05 lalpha0=-2.09415183623353e-11 alpha1=0.0 beta0=25.2626539600001 lbeta0=1.34074471872356e-5 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.3946656205 lkt1=1.52357354400379e-8 kt2=-0.019151 at=237102.9225 lat=-0.685608094801822 ute=-1.203541169 lute=2.74243237920736e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.75 nmos lmin=2e-06 lmax=4e-06 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.831727351546451+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-8.46428087113106e-9 k1=0.88325 k2=-0.0368033935204499 lk2=1.29121121475004e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=91643.7949999999 lvsat=0.0362201244004048 ua=-1.381677945785e-10 lua=-1.16991001813354e-18 ub=2.820564426195e-18 lub=-1.78489151032754e-24 uc=5.7002e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0381749445573999 lu0=-1.55022132433936e-10 a0=0.933970656530001 la0=-4.87740195175861e-7 keta=-0.020254 a1=0.0 a2=0.65972622 ags=0.16025 b0=-2.626190004485e-07 lb0=4.26734639648251e-13 b1=-7.36957729995003e-10 lb1=3.75381747273358e-15 pb1=-3.00926553810506e-36 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.04360124947+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.63455309050564e-9 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.20557 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.8066e-5 alpha1=0.0 beta0=26.388819991 lbeta0=9.04778707522128e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169000001 lkt1=6.51962239207318e-8 kt2=-0.019151 at=97424.8200000001 lat=-0.14488049760162 wat=1.11022302462516e-16 pat=-2.11758236813575e-22 ute=-1.099017662 lute=-1.30392447841457e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.76 nmos lmin=1e-06 lmax=2e-06 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.820617766536401+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.23244300926601e-8 k1=0.88325 k2=-0.0374573693387 lk2=1.41358585116182e-8 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=114920.5845 lvsat=-0.00733635846036451 ua=-1.41337023720001e-10 lua=4.76048148983641e-18 ub=1.85662102922001e-18 lub=1.88788957713363e-26 uc=5.7002e-11 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0370613347729001 lu0=1.92881015432394e-9 a0=0.282237339919998 la0=7.31809907930759e-7 keta=-0.0286126861540001 lketa=1.56411162374971e-8 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.43251245569999e-08 lb0=-1.28919381771165e-13 b1=2.10707701862e-09 lb1=-1.56805695429951e-15 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.08026278697+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.896801900253e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.73469942443 lpclm=1.75947069803982e-06 ppclm=-8.07793566946316e-28 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=2.8066e-5 alpha1=0.0 beta0=27.514255822 lbeta0=6.94182540538488e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=16515.036 lat=0.00652120752032403 ute=-1.0555257941 lute=-2.11776214222521e-7 ua1=3.0044e-9 ub1=-4.0138723e-18 lub1=4.89090564024295e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.77 nmos lmin=8.0e-07 lmax=1e-06 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.8102985436525+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=2.1314960157251e-8 k1=0.88325 k2=-0.0306811239364999 lk2=8.23211569116016e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=68433.2516489998 lvsat=0.0331653119000741 ua=-1.41632247779999e-10 lua=5.01769279509497e-18 ub=1.49004420559999e-18 lub=3.38255654158862e-25 uc=4.67991368000003e-11 luc=8.88915273723117e-18 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0406522509115002 lu0=-1.19974321318623e-9 a0=1.1222 keta=-0.0314107442740001 lketa=1.80788991920241e-8 a1=0.0 a2=0.65972622 ags=0.16025 b0=-6.05599528900001e-07 lb0=4.28609213231365e-13 b1=1.3385746724e-09 lb1=-8.9850620167645e-16 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.12712727665+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-9.9798283855821e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.8885812795 lpclm=-5.26039005732856e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.386925285e-05 lalpha0=1.23687881837128e-11 alpha1=0.0 beta0=30.52152901 lbeta0=4.32176570579874e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.379442409999999 lkt1=5.84812680081067e-9 kt2=-0.019151 at=7218.97499999986 lat=0.014620317002025 ute=-1.47144455750001 lute=1.5058926512086e-7 ua1=6.3361047035e-09 lua1=-2.90271773758206e-15 ub1=-8.9946013165e-18 lub1=4.82850589308879e-24 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.78 nmos lmin=6e-07 lmax=8.0e-07 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.783011550730507+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.96311085732052e-8 k1=0.88325 k2=-0.023096051889 lk2=3.14070434492423e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=109489.217654499 lvsat=0.00560686422257595 ua=-1.36357695470001e-10 lua=1.47719702797787e-18 ub=1.18873694125001e-18 lub=5.4050544358841e-25 uc=4.87251473850002e-11 luc=7.59633546614524e-18 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0328000283300003 lu0=4.07099052464257e-9 a0=1.1222 keta=-0.0044772 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.06056374425+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.51181118041187e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.1049 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=6.273345619e-05 lalpha0=-2.04308685304318e-11 alpha1=0.0 beta0=37.8082338000002 lbeta0=-5.6936930414571e-7 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67299999995 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210584e-8 ua1=2.0117e-9 ub1=-1.8012e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.79 nmos lmin=5e-07 lmax=6e-07 wmin=7e-07 wmax=7.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.832682109660006+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.62243047127105e-8 k1=0.88325 k2=0.00414992979899997 lk2=-9.69871931171051e-9 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=100523.184559001 lvsat=0.00983202662453175 ua=-1.68334973779999e-10 lua=1.6546201636061e-17 ub=-1.60058994799983e-19 lub=1.17611338928854e-24 uc=1.64500934039999e-10 luc=-4.69619620129438e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0390106126189997 lu0=1.1443085737099e-9 a0=1.1222 keta=0.018475888548 lketa=-1.08164364004481e-8 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.761951778700002+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=8.5600089453633e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=0.437037441000015 lpclm=3.14724220165718e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=3.76096455099999e-05 lalpha0=-8.5914988617779e-12 alpha1=0.0 beta0=35.2635323999998 lbeta0=6.2979832829164e-7 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.444978200000001 lkt1=3.49887960161979e-8 kt2=-0.019151 at=29133.8246399998 lat=0.00436660174282189 ute=-1.879349683 lute=2.73437440866603e-7 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=-1.06577157899999e-18 lub1=-3.4656402454046e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.80 nmos lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.838095495661428+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' wvth0=-5.23770517643172e-9 k1=0.88325 k2=-0.0350098659205714 wk2=9.44035163456431e-10 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=68129.2014285714 wvsat=0.0201257380997314 ua=-3.20773584885714e-10 wua=1.11618651310806e-16 ub=2.82081495784286e-18 wub=-2.8244838660853e-25 uc=3.19430594428571e-11 wuc=1.53427874170407e-17 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0373452888314285 wu0=4.83453650958896e-10 a0=0.456701523714286 wa0=2.15076570118502e-7 keta=-0.0266193055428571 wketa=3.89727289411406e-9 a1=0.0 a2=0.65972622 ags=0.16025 b0=-3.31415371742857e-07 wb0=1.09613343110256e-13 b1=8.78174185714286e-11 wb1=8.87130910461085e-17 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.855558035428571+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' wnfactor=1.1665662488422e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.143786068571429 wpclm=2.13899541392091e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=1.69635021142857e-05 walpha0=6.79770417549051e-12 alpha1=0.0 beta0=34.0161812285714 wbeta0=-3.23900868045497e-6 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.394290014285714 wkt1=2.17968282668573e-9 kt2=-0.019151 at=-177334.285714286 wat=0.145312188445714 ute=-1.24400978 wute=6.81514163810401e-8 ua1=3.0044e-9 ub1=-4.10873876285714e-18 wub1=2.18113594857017e-25 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.81 nmos lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.876877861632547+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-7.70653740762307e-07 wvth0=-1.92190269829696e-08 pvth0=2.77826215116273e-13 k1=0.88325 k2=-0.0308621305233539 lk2=-8.24206496823391e-08 wk2=-6.11146632625018e-10 pk2=3.09033922687473e-14 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=52495.1335916639 lvsat=0.310668329797538 wvsat=0.025320438551765 pvsat=-1.03225144605168e-7 ua=-3.0908883758901e-10 lua=-2.32190429556901e-16 wua=1.07046600045982e-16 pua=9.08523325476775e-23 ub=3.93536677584284e-18 lub=-2.21475277824657e-23 wub=-7.33642434485312e-25 pub=8.96578566312506e-30 uc=3.81909493050195e-11 luc=-1.24153325192484e-16 wuc=1.32668135483198e-17 puc=4.12521770550562e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0391269077420172 lu0=-3.54029787424637e-08 wu0=-2.20785693809002e-10 pu0=1.39941097415649e-14 a0=-0.144844855610945 la0=1.19534730762491e-05 wa0=4.58335670909411e-07 pa0=-4.83386021725945e-12 keta=-0.0243473455929799 lketa=-4.51466637063577e-08 wketa=3.14237330548826e-09 pketa=1.5000791656384e-14 a1=0.0 a2=0.65972622 ags=0.144258786943699 lags=3.17765248524106e-07 wags=5.31336837979105e-09 pags=-1.05583223596607e-13 b0=-5.85096029118562e-07 lb0=5.04094947975105e-12 wb0=1.90507696755043e-13 pb0=-1.60747119681479e-18 b1=1.7045958733931e-09 lb1=-3.21273943193691e-14 wb1=-8.07730170447026e-16 pb1=1.78134400919561e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.80125414652002+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.07908566373905e-06 wnfactor=1.46752527044396e-07 pnfactor=-5.98042924937283e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.32312548118982 lpclm=2.34349376889385e-05 wpclm=6.05756289343979e-07 ppclm=-7.78667987602821e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=7.45220717440168e-08 lalpha0=3.35604992669536e-10 walpha0=1.60342628416247e-11 palpha0=-1.83541883265391e-16 alpha1=0.0 beta0=37.3275247684563 lbeta0=-6.58005055148463e-05 wbeta0=-4.55960638252699e-06 pbeta0=2.62419152019194e-11 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.403097098987989 lkt1=1.7500770262632e-07 wkt1=8.3751971272762e-09 pkt1=-1.2311255778598e-13 kt2=-0.019151 at=-359352.854441936 lat=3.6169348456622 wat=0.220611516099045 pat=-1.4962910869373e-6 ute=-1.25301023766733 lute=1.78850263417857e-07 wute=8.81200355498663e-08 pute=-3.96801243940968e-13 ua1=3.0044e-9 ub1=-4.34240885918968e-18 lub1=4.64331479871702e-24 wub1=3.61182317398346e-25 pub1=-2.84295306518087e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.82 nmos lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.737552072173816+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=3.26013125582632e-07 wvth0=2.7030176109881e-08 pvth0=-8.62124084854983e-14 k1=0.88325 k2=-0.0441931551184891 lk2=2.25110576828968e-08 wk2=3.61363769378075e-09 pk2=-2.35090333741528e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=108140.568307572 lvsat=-0.127330297401145 wvsat=0.00876067550646151 pvsat=2.71207412273096e-8 ua=-3.53774357459573e-10 lua=1.19540066554585e-16 wua=1.24077531553956e-16 pua=-4.32022338060746e-23 ub=-2.82985403152891e-19 lub=1.10561388412848e-23 wub=9.24278158938325e-25 pub=-4.0841068865754e-30 uc=-1.50679704797229e-11 luc=2.95060467832892e-16 wuc=3.88779092014627e-17 puc=-1.60338929104884e-22 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0330611615518391 lu0=1.23419713652601e-08 wu0=1.94672098503749e-09 pu0=-3.06685769674536e-15 a0=2.0327256717049 la0=-5.18670933875101e-06 wa0=-3.74727089566043e-07 pa0=1.72337753856812e-12 keta=-0.0400848427420999 lketa=7.87269690911784e-08 wketa=1.02333440661232e-08 pketa=-4.08139481245267e-14 a1=0.0 a2=0.65972622 ags=0.208223639168903 lags=-1.85717518869864e-07 wags=-1.59401051393731e-08 pags=6.17079885598519e-14 b0=4.16528268420126e-07 lb0=-2.84307675763166e-12 wb0=-1.25050028309092e-13 pb0=8.76359706576748e-19 b1=-4.23329020784967e-09 lb1=1.46111380566383e-14 wb1=2.45401366680883e-15 pb1=-7.86053173134955e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.936859226979205+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.17053946204179e-08 wnfactor=7.63364008181501e-08 pnfactor=-4.37806251240856e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=3.39423216928374 lpclm=-1.36965212611327e-05 wpclm=-9.6167070246357e-07 ppclm=4.55091572639403e-12 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.14670840240364e-05 lalpha0=9.79416193561188e-12 walpha0=-4.89298481357064e-12 palpha0=-1.88184735046638e-17 alpha1=0.0 beta0=26.4525984102288 lbeta0=1.97986607080147e-05 wbeta0=-7.28564908652704e-07 pbeta0=-3.9131355199404e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37131417849475 lkt1=-7.51633242598054e-08 wkt1=-1.42973406936703e-08 pkt1=5.5348451484305e-14 kt2=-0.019151 at=161996.321517022 lat=-0.486730163462161 wat=0.0459853683706463 pat=-1.21766593265472e-7 ute=-1.32473515300725 lute=7.43414357762931e-07 wute=7.42031982001495e-08 pute=-2.87258463203545e-13 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.83 nmos lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.818199639991855+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=1.38069544951579e-08 wvth0=8.28258489810874e-09 pvth0=-1.36359647352468e-14 k1=0.88325 k2=-0.0389878796044437 lk2=2.36018169662816e-09 wk2=1.33749092567463e-09 pk2=6.4606093532946e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=52569.7356159714 lvsat=0.0877977885187213 wvsat=0.0239237961909404 pvsat=-3.15793532543932e-8 ua=-3.99539585267726e-10 lua=2.96708292819849e-16 wua=1.60029583541711e-16 pua=-1.82381291495205e-22 ub=3.38481551745301e-18 lub=-3.14280246240253e-24 wub=-3.45472887142361e-25 pub=8.31405422805036e-31 uc=6.92511632597751e-11 luc=-3.13592197839362e-17 wuc=-7.49977069073598e-18 puc=1.92002467786711e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.03557330788042 lu0=2.61684750005808e-09 wu0=1.59289888494119e-09 pu0=-1.69712707614651e-15 a0=0.860768328963871 la0=-6.49780023280897e-07 wa0=4.48194426942587e-08 pa0=9.9211801474219e-14 keta=-0.0197484779714286 wketa=-3.09514961389371e-10 a1=0.0 a2=0.65972622 ags=0.16025 b0=-5.75993014518294e-07 lb0=9.99212326252149e-13 wb0=1.91868880846485e-13 pb0=-3.50509768221595e-19 b1=-2.13282731911063e-09 lb1=6.47974000277335e-15 wb1=8.54646281588652e-16 pb1=-1.66899513562239e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.893027602964041+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.813881746045e-07 wnfactor=9.219142539891e-08 pnfactor=-1.0515924633713e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.143786068571428 wpclm=2.13899541392091e-7 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.54104428773938e-05 lalpha0=-5.47153053521804e-12 walpha0=-1.06194473516561e-11 palpha0=3.35004305773689e-18 alpha1=0.0 beta0=30.4432409990619 lbeta0=4.34992150177789e-06 wbeta0=-2.48239224176406e-06 pbeta0=2.87635275892098e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.407571169 lkt1=6.51962239207292e-8 kt2=-0.019151 at=51485.9091218571 lat=-0.0589177240710931 wat=0.0281269250855388 pat=-5.26322554239887e-8 ute=-1.099017662 lute=-1.30392447841458e-7 ua1=3.0044e-9 ub1=-3.7525e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.84 nmos lmin=1e-06 lmax=2e-06 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.825665272606629+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-1.63043344544095e-10 wvth0=-3.09042644660725e-09 pvth0=7.6456803864503e-15 k1=0.88325 k2=-0.0454197063875077 lk2=1.43956796779958e-08 wk2=4.87508418019942e-09 pk2=-1.59080185895588e-16 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=111215.641498712 lvsat=-0.0219428350512044 wvsat=0.00226841804151248 pvsat=8.94307820932044e-9 ua=-2.43601942824849e-10 lua=4.91138283739765e-18 wua=6.2613537490488e-17 pua=-9.23920662684959e-26 ub=1.57103984962724e-18 lub=2.51208932035441e-25 wub=1.748522176669e-25 pub=-1.42248246643349e-31 uc=5.24926485714286e-11 wuc=2.76093158046857e-18 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0364445996674886 lu0=9.86450585132052e-10 wu0=3.77607169520021e-10 pu0=5.76976608709912e-16 a0=-0.0167816848222144 la0=9.92327542066191e-07 wa0=1.83079780240866e-07 pa0=-1.59506610816833e-13 keta=-0.027666732607734 lketa=1.48169627238948e-08 wketa=-5.79177085865207e-10 pketa=5.04602823466289e-16 a1=0.0 a2=0.65972622 ags=0.16025 b0=1.21866075426608e-07 lb0=-3.06650215075441e-13 wb0=-5.35985229070334e-14 pb0=1.08818901845543e-19 b1=6.62625748645737e-09 lb1=-9.91061860788254e-15 wb1=-2.76694958668185e-15 pb1=5.10788353851598e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.08645424141056+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.80559681748793e-07 wnfactor=-3.79082942741087e-09 pnfactor=7.44466841663295e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-1.54195952865152 lpclm=2.61631950361373e-06 wpclm=4.94259529491501e-07 ppclm=-5.24621104491127e-13 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=4.09904114673613e-05 lalpha0=2.79941346052257e-12 walpha0=-7.91320356029836e-12 palpha0=-1.71399128064723e-18 alpha1=0.0 beta0=27.3460153662938 lbeta0=1.01455770920645e-05 wbeta0=1.03008247334302e-07 pbeta0=-1.96155463769995e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37273 kt2=-0.019151 at=16515.036 lat=0.00652120752032401 ute=-1.0555257941 lute=-2.11776214222522e-7 ua1=3.0044e-9 ub1=-4.32403534063e-18 lub1=1.06948036233582e-24 wub1=1.89902904560449e-25 pub1=-3.55354101032599e-31 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.81e-6 sbref=2.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.85 nmos lmin=8.0e-07 lmax=1e-06 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.755518949506103+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=6.09513093398815e-08 wvth0=3.35397925488262e-08 pvth0=-2.42680682413503e-14 k1=0.88325 k2=-0.0288349219835414 lk2=-5.36644709002979e-11 wk2=-1.1303703773341e-09 pk2=5.07311804826446e-15 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=15923.8398695603 lvsat=0.0610792894919794 wvsat=0.0321498325313739 pvsat=-1.7090835232241e-8 ua=-4.2130236482708e-10 lua=1.59731276203043e-16 wua=1.71233063224182e-16 pua=-9.47261762860178e-23 ub=2.29515189622959e-18 lub=-3.7966717155844e-25 wub=-4.929416755264e-25 pub=4.39561172656275e-31 uc=-3.71851037501013e-12 luc=4.89734663316543e-17 wuc=3.09303388005492e-17 puc=-2.45423425158302e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0315018332508821 lu0=5.29279134070273e-09 wu0=5.60250792023124e-09 pu0=-3.97517114624045e-15 a0=1.1222 keta=-0.0560350596255479 lketa=3.9532612323222e-08 wketa=1.50766803116616e-08 pketa=-1.31354220314123e-14 a1=0.0 a2=0.65972622 ags=0.16025 b0=-1.11290736753844e-06 lb0=7.69135034146869e-13 wb0=3.10608355747479e-13 pb0=-2.08493063320294e-19 b1=-2.06877570456196e-08 lb1=1.38864707270588e-14 wb1=1.34860180683284e-14 pb1=-9.05236825420285e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='1.04326239218623+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.42929171838741e-07 wnfactor=5.1347785080864e-08 pnfactor=2.64076625235253e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=2.78129198013181 lpclm=-1.15027446415017e-06 wpclm=-5.46578195254434e-07 ppclm=3.82199395654246e-13 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=-5.27764624119503e-06 lalpha0=4.31100423265829e-11 walpha0=1.17230336127678e-11 palpha0=-1.88218861915466e-17 alpha1=0.0 beta0=28.1440672281953 lbeta0=9.45028158984962e-06 wbeta0=1.45564377022202e-06 pbeta0=-3.14002616329616e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37944241 lkt1=5.84812680081025e-9 kt2=-0.019151 at=7218.97500000001 lat=0.014620317002025 ute=-1.4714445575 lute=1.50589265120858e-7 ua1=6.3361047035e-09 lua1=-2.90271773758205e-15 ub1=-7.44378611335e-18 lub1=3.78753514531117e-24 wub1=-9.49514522802244e-25 pub1=6.373530778003e-31 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.41e-6 sbref=2.41e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.86 nmos lmin=6e-07 lmax=8.0e-07 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.768341210028917+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=5.2344482364287e-08 wvth0=8.98218016067705e-09 pvth0=-7.78399194431609e-15 k1=0.88325 k2=-0.0319918861567214 lk2=2.06541931766923e-09 wk2=5.44663465542922e-09 pk2=6.58362613067379e-16 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=68859.7320644314 lvsat=0.0255465482792019 wvsat=0.02487613388326 pvsat=-1.22084304779824e-8 ua=-1.68278135973694e-10 lua=-1.01089601967323e-17 wua=1.95438642663161e-17 pua=7.09383331165908e-24 ub=-4.35052247420504e-19 lub=1.45295778802939e-24 wub=9.94194158968911e-25 pub=-5.58665372026192e-31 uc=4.44948386397113e-11 luc=1.66106897256636e-17 wuc=2.59008267486038e-18 puc=-5.51920065376678e-24 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.029896894678566 lu0=6.37009191292272e-09 wu0=1.77749583449616e-09 pu0=-1.40766620879957e-15 a0=1.1222 keta=0.00285975210857144 wketa=-4.49218099361081e-9 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.823808911974293+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.3770016721988e-09 wnfactor=1.44957407647782e-07 pnfactor=-3.64269541379148e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=2.27496908716247 lpclm=-8.10409779150537e-07 wpclm=-7.16395859858793e-07 ppclm=4.96187974660941e-13 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=0.000125503457420496 lalpha0=-4.46755964763944e-11 walpha0=-3.84320631133934e-11 palpha0=1.48442710900186e-17 alpha1=0.0 beta0=47.7153459414405 lbeta0=-3.68676310490783e-06 wbeta0=-6.0658077366155e-06 pbeta0=1.90868046760496e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.37073 kt2=-0.019151 at=6851.67299999998 lat=0.014866865163807 ute=-1.12457734 lute=-8.22422328210592e-8 ua1=2.0117e-9 ub1=-1.8012e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=2.02e-6 sbref=2.01e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__nfet_g5v0d10v5__model.87 nmos lmin=5e-07 lmax=6e-07 wmin=4.2e-07 wmax=7.0e-7 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=6.43795e-8 ll=0.0 lw=0.0 lwl=0.0 wint=4.3866e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.20872e-08+sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre*(1.20872e-08*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='0.87993839021345+sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))' lvth0=-2.44684423051775e-10 wvth0=-2.89335083818999e-08 pvth0=1.0083435040176e-14 k1=0.88325 k2=-0.00898356822880039 lk2=-8.77704343100219e-09 wk2=8.0412205704853e-09 pk2=-5.64312648129555e-16 k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90875.2361210983 lvsat=0.0151719401320342 wvsat=0.00590713009417726 pvsat=-3.26945816341118e-9 ua=-5.06651181788546e-10 lua=1.49346292286104e-16 wua=2.07140188044977e-16 pua=-8.13092459021208e-23 ub=1.19752281510754e-18 lub=6.83621482988614e-25 wub=-8.3120389958847e-25 pub=3.01537034486447e-31 uc=2.34709527400798e-10 luc=-7.30262704207996e-17 wuc=-4.29864750398289e-17 puc=1.59583419802611e-23 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.0486596465479778 lu0=-2.47168604077074e-09 wu0=-5.90779470562738e-09 pu0=2.21395779061879e-15 a0=1.1222 keta=0.053050615033953 lketa=-2.36519924358198e-08 wketa=-2.11689986361015e-08 pketa=7.85880022266496e-15 a1=0.0 a2=0.65972622 ags=0.16025 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))' nfactor='0.402411058330014+sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.02956947621383e-07 wnfactor=2.20135277779491e-07 pnfactor=-7.1853848836652e-14 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-8.0e-4 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.032 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=-0.228931611897256 lpclm=3.69530890175069e-07 wpclm=4.07751540079297e-07 ppclm=-3.35563702332851e-14 pdiblc1=0.21098 pdiblc2=2.0e-4 pdiblcb=-0.26831 drout=0.36075 pscbe1=937310000.0 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=9.09603475489768e-05 lalpha0=-2.83974668374297e-11 walpha0=-3.26649276360003e-11 palpha0=1.21265604005164e-17 alpha1=0.0 beta0=50.7759687188254 lbeta0=-5.12905404314546e-06 wbeta0=-9.4977683600546e-06 pbeta0=3.52596102375503e-12 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.378897036827857 lkt1=3.8486426017965e-09 wkt1=-4.04593816130816e-08 pkt1=1.90661194507301e-14 kt2=-0.019151 at=67478.5209233554 lat=-0.0137029912784429 wat=-0.0234772305040174 pat=1.10634335799437e-8 ute=-2.56571269781465 lute=5.96879834330877e-07 wute=4.20238110354539e-07 pute=-1.98033427361584e-13 ua1=-1.673609407e-09 lua1=1.73666889026409e-15 ub1=-8.78933793056004e-18 lub1=3.29309710653505e-24 wub1=4.72889252293697e-24 pub1=-2.22844804140134e-30 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo=3.059976892e-10 cgso=3.059976892e-10 cgbo=0.0 capmod=2.0 xpart=0.0 cgsl=4.9879e-11 cgdl=4.9879e-11 cf=0.0 clc=1.0e-7 cle=0.6 dlc=5.38675e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.00095274816 mjs=0.295 pbs=0.72468 cjsws=1.005492404e-10 mjsws=0.037586 pbsws=0.29067 cjswgs=6.37254e-11 mjswgs=0.78692 pbswgs=0.54958 saref=1.81e-6 sbref=1.81e-6 wlod='0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff' kvth0='0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff' lkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff' wkvth0='0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff' lku0='0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff' wku0='0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff' steta0=0.0 tku0=0.0
.ends sky130_fd_pr__nfet_g5v0d10v5