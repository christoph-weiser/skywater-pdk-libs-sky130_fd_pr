* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b=-0.029
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=1.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=1.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=0.89805
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=9.9505e-1
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=1.0144
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_0='-0.015262+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_0=-3503.4
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_0=0.0013127
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_0=-0.0029685
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_1='-0.0025365+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_1=323.35
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_1=-0.00053421
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_1=-0.0010115
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_0=-3946.4
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_0='-0.024526+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_0=0.0010173
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_0=-0.0031271
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_1=-1841.7
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_1='-0.0099998+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_1=-0.00057848
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_1=-0.0013993
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_2=-2994.9
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_2='-0.0082165+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_2=-0.0015137
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_2=-0.003002
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_0=0.00059498
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_0=-0.0016449
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_0='-0.015075+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_0=1100.9
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_1=-0.0068059
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_1=-0.002939
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_1='-0.012671+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_1=-3862.9
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_2=-0.0017173
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_2=-0.0041054
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_2='-0.022123+sky130_fd_pr__nfet_g5v0d10v5__vth0_correldiff_rf_b'
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_2=-5556.8
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"