* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope=2.0e-3
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope=0.0255
.param sky130_fd_bs_flash__special_sonosfet_star__tox_slope1=2.0e-3
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_slope1=0.028