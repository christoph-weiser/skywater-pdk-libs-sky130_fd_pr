* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__ind_03_90 a b ct sub
r31 net27 b r='1e-2'
r26 a net23 r='1e-2'
c24 net35 net27 c='8.337e-15'
c25 net23 net37 c='53.8e-15'
c0 net27 net31 c='53.8e-15'
r1 sub net31 r='21.56'
r13 net23 net35 r='50.11'
r10 sub net37 r='21.56'
r0 net41 net27 r='1.019'
r9 net23 net39 r='1.019'
l0 ct net41 l=760.5e-12
l1 net39 ct l=760.5e-12
.ends sky130_fd_pr__ind_03_90