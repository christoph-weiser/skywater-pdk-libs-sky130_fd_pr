* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff=-0.034
.param sky130_fd_pr__nfet_05v0_nvt__toxe_mult=1.0
.param sky130_fd_pr__nfet_05v0_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_05v0_nvt__overlap_mult=7.7117e-1
.param sky130_fd_pr__nfet_05v0_nvt__ajunction_mult=9.7602e-1
.param sky130_fd_pr__nfet_05v0_nvt__pjunction_mult=1.0437e+0
.param sky130_fd_pr__nfet_05v0_nvt__lint_diff=0.0
.param sky130_fd_pr__nfet_05v0_nvt__wint_diff=0.0
.param sky130_fd_pr__nfet_05v0_nvt__dlc_diff=-1.5781e-8
.param sky130_fd_pr__nfet_05v0_nvt__dwc_diff=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0=0.010308
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_0=0.0064317
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_0=-0.00025708
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_0=-0.0078378
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_0=-2.691e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0='-0.0046033+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_0=0.00034013
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_0=-1.3689e-18
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_1=-1.2472e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1=0.029952
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_1=-0.00044213
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_1=-0.0039719
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_1=-0.0070434
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_1=-2.4351e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1='-0.0022002+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_1=-0.00056708
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_2=-1.5224e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2=-0.044586
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_2=0.0015915
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_2=-0.008363
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_2=-3.3419e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2=-2848.5
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2='-0.0011931+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_3=-1.6915e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_3=0.0075894
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_3=-9.6861e-19
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3=0.064023
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_3=0.0012767
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_3=-0.0046305
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_3=-0.0066322
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3='-0.013446+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_4=-0.0078468
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4='-0.0057166+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_4=-2.429e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_4=-0.0084686
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_4=-1.2894e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4=0.024393
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_4=-0.035687
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_4=-0.0016893
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_5=-0.00013553
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_5=-0.0079399
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5='-0.0050535+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_5=-2.1501e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_5=0.0053237
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_5=-1.2037e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5=0.053081
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_5=0.02762
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_6=0.00043703
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_6=-0.0023615
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_6=-0.0068188
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6='-0.011078+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_6=-1.9014e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_6=-0.00041719
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_6=-1.0585e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6=0.055346
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7=0.0016268
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_7=0.00035232
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_7=-0.0094947
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7='-0.014254+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_7=-2.898e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7=-3146.5
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_7=-1.429e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8=0.017467
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_8=8.0096e-8
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_8=-0.0049283
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_8=-0.0086023
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8='-0.031553+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_8=-2.2873e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_8=1.6514e-9
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_8=-1.2296e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9=-0.011611
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_9=-0.0030036
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_9=-0.0089225
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9='-0.010333+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_9=-1.3766e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9=-6052.7
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_9=-9.127e-19
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10=-4889.9
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10='-0.010495+sky130_fd_pr__nfet_05v0_nvt__vth0_correldiff'
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10=0.011275
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_10=-0.0096426
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_10=0.00063457
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_10=-2.505e-11
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_10=-1.3111e-18
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10=0.0
.include "sky130_fd_pr__nfet_05v0_nvt.pm3.spice"