* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult=0.948
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult=0.8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult=0.86067
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult=0.82447
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult=0.75
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff=1.7325e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff=-3.2175e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff=-7.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff=-6.425e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff=1.1336e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42=0.85
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42=0.65
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42=0.65
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult=0.85
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult=0.75
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult=0.75
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_0=-0.065542
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_0=0.0010442
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_0=-32505.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_0=-0.21576
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_0=-2.0987
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_0=-0.0038838
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_1=-0.28484
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_1=-0.21491
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_1=0.0043607
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_1=-0.059034
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_1=0.00085042
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_1=-26494.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_2=-0.13248
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_2=0.047598
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_2=-0.0034116
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_2=-0.042789
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_2=0.0016287
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_2=-20516.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_3=-0.17311
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_3=-1.9691
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_3=0.016626
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_3=-0.073889
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_3=-0.0038
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_3=-37673.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_4=-0.31537
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_4=0.4484
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_4=0.010615
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_4=-0.067217
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_4=-0.0036293
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_4=-25995.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_5=-0.079709
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_5=0.96083
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_5=0.0050505
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_5=-0.029865
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_5=-0.00025925
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_5=-18682.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_6=-0.047966
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_6=-1.5615
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_6=0.0032612
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_6=-0.064411
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_6=-0.0093565
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_6=-31246.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_7=-0.15151
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_7=0.22325
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_7=0.0089861
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_7=-0.056878
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_7=-0.0052178
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_7=-22366.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_8=-0.20897
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_8=1.5448
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_8=0.0046298
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_8=-0.02487
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_8=-0.00059818
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_8=-16469.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_0=-2.2103
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_0=-0.0043971
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_0=-0.068994
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_0=-0.0051783
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_0=-28908.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_0=-0.21764
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_1=0.038663
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_1=0.0032931
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_1=-0.066959
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_1=-0.0030718
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_1=-26301.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_1=-0.24936
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_2=0.37546
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_2=0.0033757
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_2=-0.048089
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_2=-0.00068406
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_2=-15222.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_2=-0.10997
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_3=-0.15284
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_3=-1.8412
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_3=0.014866
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_3=-0.072281
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_3=-0.0047778
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_3=-38008.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_4=-0.008134
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_4=-24439.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_4=-0.26445
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_4=-0.60655
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_4=0.0080453
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_4=-0.062068
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_5=-0.041218
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_5=-0.0034389
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_5=-9878.8
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_5=-0.091057
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_5=1.0698
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_5=0.0034441
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_6=0.0075537
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_6=-0.069722
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_6=-0.0070527
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_6=-35711.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_6=0.0093774
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_6=-2.2074
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_7=0.80674
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_7=0.0046426
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_7=-0.055588
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_7=-0.0090538
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_7=-24756.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_7=-0.12664
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_8=1.1546
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_8=0.0027331
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_8=-0.005212
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_8=-7446.5
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_8=-0.041012
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_8=-0.18505
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_8=0.0
.include "sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"