* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre=0.0
.subckt sky130_fd_pr__pfet_01v8_lvt d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-0.54483+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' k1=0.64774 k2=-0.075662 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.0054e-9 ub=3.0419e-18 uc=4.9353e-11 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=0.00266747 a0=1.75814 keta=-0.01258 a1=0.0 a2=0.46703705 ags=0.412557 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=0.0018466 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=0.01363 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.60135 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-0.54483+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' k1=0.64774 k2=-0.075662 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.0054e-9 ub=3.0419e-18 uc=4.9353e-11 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=0.00266747 a0=1.75814 keta=-0.01258 a1=0.0 a2=0.46703705 ags=0.412557 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=0.0018466 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=0.01363 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.60135 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.569562915e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=9.723654767e-8 k1=0.64774 k2=-7.570419588e-02 lk2=3.383541841e-10 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.064574695e-09 lua=4.745014629e-16 ub=3.131516007e-18 lub=-7.185998386e-25 uc=3.772200777e-11 luc=9.326491403e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.582405120e-03 lu0=6.821059230e-10 a0=1.842411195e+00 la0=-6.757416419e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.987800460e-01 lags=1.104726411e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=6.412557475e-05 lpdiblc2=1.429304746e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.812711361e-03 ldelta=6.268414063e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.113966375e-01 lkt1=8.056052002e-8 kt2=-0.055045 at=2.992533804e+05 lat=-1.094817467e-1 ute=-3.128584783e-01 lute=7.228695462e-7 ua1=6.681850806e-10 lua1=1.121402439e-16 ub1=-1.755248019e-19 lub1=2.155799516e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.197901416e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.212138621e-8 k1=0.64774 k2=-5.288086075e-02 lk2=-9.138075563e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.570799194e+05 lvsat=-1.339012608e-1 ua=-3.115158625e-09 lua=6.777808277e-16 ub=3.178587495e-18 lub=-9.077639092e-25 uc=6.137107612e-11 luc=-1.772532745e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.486071178e-03 lu0=1.069238803e-9 a0=2.303320336e+00 la0=-2.527976466e-6 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.416218713e-01 lags=-6.169387426e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.229999040e-04 lpdiblc2=1.365458634e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.965880746e-02 ldelta=7.041457312e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.59135 kt2=-0.055045 at=3.793216998e+05 lat=-4.312486990e-1 ute=-0.13298 ua1=6.9609e-10 ub1=-1.575546805e-19 lub1=1.433642331e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos lmin=1.5e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.554205113e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.980403769e-8 k1=0.64774 k2=-1.461324234e-01 lk2=9.686197752e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90748.0 ua=-2.226002118e-09 lua=-1.117119401e-15 ub=1.817403269e-18 lub=1.839997434e-24 uc=2.695198567e-11 luc=6.770773628e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.238075017e-03 lu0=-4.487975080e-10 a0=1.152012669e+00 la0=-2.038834877e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.460547025e-01 lags=5.349542688e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-3.445352388e-03 lpdiblc2=2.105972404e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.686888023e-02 ldelta=1.267335786e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.59135 kt2=-0.055045 at=2.064810733e+05 lat=-8.234310407e-2 ute=-0.13298 ua1=8.017883880e-10 lua1=-2.133685794e-16 ub1=-3.161404494e-19 lub1=4.634941886e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos lmin=1e-06 lmax=1.5e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.330898664e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.410850784e-8 k1=0.64774 k2=-5.135944028e-02 lk2=-4.706548713e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=9.000845647e+04 lvsat=1.123111480e-3 ua=-3.157792953e-09 lua=2.979494090e-16 ub=3.143700553e-18 lub=-1.741905683e-25 uc=6.931940672e-11 luc=3.366240468e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.143048399e-03 lu0=1.214170141e-9 a0=8.322710737e-01 la0=2.816936853e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-9.515840300e-02 lags=9.012737576e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.522571395e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.501727831e-8 nfactor='2.599234224e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-9.405671895e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=3.576886000e-04 lpdiblc2=1.528421683e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=9.871018390e-03 ldelta=2.330069574e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.524693000e-01 lkt1=9.281913054e-8 kt2=-9.429581446e-02 lkt2=5.960844563e-8 at=2.056171489e+05 lat=-8.103110096e-2 ute=6.076818100e-02 lute=-2.942366438e-7 ua1=6.6129e-10 ub1=-1.049382911e-20 lub1=-6.775796530e-28 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos lmin=5e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.596055551e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.290183103e-8 k1=0.64774 k2=-1.186069080e-01 lk2=2.143648207e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=4.236987772e+04 lvsat=4.965038792e-2 ua=-2.786153247e-09 lua=-8.062323568e-17 ub=2.817829617e-18 lub=1.577594900e-25 uc=7.591434732e-11 luc=-3.351728749e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.404884209e-03 lu0=-7.120521602e-11 a0=1.179367975e+00 la0=-7.187830909e-8 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.172107689e+00 lags=-3.896331838e-7 b0=1.380555879e-06 lb0=-1.406310149e-12 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.115428605e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=1.537441781e-8 nfactor='2.475365776e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.212249495e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-2.461696471e-02 lpdiblc2=4.072477230e-08 ppdiblc2=-2.524354897e-29 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.081074845e-02 ldelta=1.215688501e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-4.881055409e-01 lkt1=-7.461083448e-8 kt2=-1.478799484e-02 lkt2=-2.138259236e-8 at=1.952938455e+05 lat=-7.051521638e-2 ute=-5.132237600e-02 lute=-1.800550375e-7 ua1=4.174599114e-10 lua1=2.483787389e-16 ub1=5.988425559e-19 lub1=-6.213811349e-25 wub1=2.295887404e-40 pub1=-2.299005293e-46 uc1=-2.348171346e-11 luc1=1.377294237e-17 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos lmin=3.5e-07 lmax=5e-07 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.495253540e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=7.673684329e-9 k1=0.64774 k2=-8.591481550e-02 lk2=4.480564853e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=2.142115113e+05 lvsat=-3.947613455e-2 ua=-3.083409290e-09 lua=7.355009730e-17 ub=3.023692000e-18 lub=5.098793574e-26 uc=8.496991780e-11 luc=-8.048445657e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.430105233e-03 lu0=4.343687740e-10 a0=1.141011921e+00 la0=-5.198474988e-8 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.104247750e-01 lags=5.417468172e-9 b0=-4.601852930e-06 lb0=1.696496092e-12 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-9.851618090e-02 lpdiblc2=7.905297027e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.353404670e-02 ldelta=1.074443276e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.565370000e-01 lkt1=1.274698394e-8 kt2=-0.056015 at=1.431951817e+05 lat=-4.349398388e-02 wat=2.220446049e-16 ute=-0.39848 ua1=8.9635e-10 ub1=-5.9922e-19 uc1=3.0734e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.897593728e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=3.118102064e-7 k1=0.64774 k2=-8.192840015e-02 wk2=4.348886716e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.120749187e-09 wua=8.005242792e-16 ub=3.230361305e-18 wub=-1.307922966e-24 uc=5.085723244e-11 wuc=-1.043938514e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.776145236e-03 wu0=-7.542070072e-10 a0=1.739392670e+00 wa0=1.301066227e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.849207072e-01 wags=-5.022047068e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.346281809e-03 wpdiblc2=-3.467795753e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.577083720e-03 wdelta=6.976731941e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.60135 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.897593728e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=3.118102064e-7 k1=0.64774 k2=-8.192840015e-02 wk2=4.348886716e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.120749187e-09 wua=8.005242792e-16 ub=3.230361305e-18 wub=-1.307922966e-24 uc=5.085723244e-11 wuc=-1.043938514e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.776145236e-03 wu0=-7.542070072e-10 a0=1.739392670e+00 wa0=1.301066227e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.849207072e-01 wags=-5.022047068e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.346281809e-03 wpdiblc2=-3.467795753e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.577083720e-03 wdelta=6.976731941e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.60135 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-6.233508423e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.693584055e-07 wvth0=4.607787142e-07 pvth0=-1.194527070e-12 k1=0.64774 k2=-9.954970837e-02 lk2=1.412991912e-07 wk2=1.654880474e-07 pk2=-9.782693369e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.326085615e-09 lua=1.646521974e-15 wua=1.814887876e-15 pua=-8.133831726e-21 ub=3.541329206e-18 lub=-2.493544314e-24 wub=-2.844106885e-24 pub=1.231812886e-29 uc=1.049764286e-11 luc=3.236296247e-16 wuc=1.889373102e-16 puc=-1.598732935e-21 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.561276826e-03 lu0=1.722955650e-09 wu0=1.466305312e-10 pu0=-7.223505431e-15 a0=2.045313542e+00 la0=-2.453073935e-06 wa0=-1.408143911e-06 pa0=1.233470034e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.561533031e-01 lags=-5.711896112e-07 wags=-1.092171663e-06 pags=4.730741484e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.402008277e-04 lpdiblc2=1.993824643e-08 wpdiblc2=1.418026867e-09 ppdiblc2=-3.917772599e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-1.186344505e-02 ldelta=1.238122732e-07 wdelta=1.226726669e-07 pdelta=-4.242297294e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.113966375e-01 lkt1=8.056052002e-8 kt2=-0.055045 at=2.992533804e+05 lat=-1.094817467e-1 ute=-3.128584783e-01 lute=7.228695462e-7 ua1=6.681850806e-10 lua1=1.121402439e-16 ub1=-1.755248020e-19 lub1=2.155799516e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.483649961e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.198384028e-08 wvth0=1.983097189e-07 pvth0=-1.397547298e-13 k1=0.64774 k2=1.404482721e-02 lk2=-3.151980571e-07 wk2=-4.644648099e-07 pk2=1.553293863e-12 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=2.393802537e+05 lvsat=-4.646379106e-01 wvsat=-5.711649782e-01 pvsat=2.295314996e-6 ua=-3.649200199e-09 lua=2.945008013e-15 wua=3.706252793e-15 pua=-1.573457481e-20 ub=4.000342353e-18 lub=-4.338159793e-24 wub=-5.702985293e-24 pub=2.380697487e-29 uc=1.107891348e-10 luc=-7.940728070e-17 wuc=-3.429617224e-16 puc=5.387857719e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.322756937e-03 lu0=2.681484793e-09 wu0=1.133402135e-09 pu0=-1.118900007e-14 a0=3.559720686e+00 la0=-8.538953776e-06 wa0=-8.719428479e-06 pa0=4.171623062e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=8.709134905e-01 lags=-1.836102212e-06 wags=-2.979287272e-06 pags=1.231440806e-11 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.326152705e-03 lpdiblc2=1.002682247e-08 wpdiblc2=-1.459589726e-08 ppdiblc2=2.517671029e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.351569574e-02 ldelta=-5.855083780e-08 wdelta=-9.616691553e-08 pdelta=4.552110528e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.59135 kt2=-0.055045 at=5.833523358e+05 lat=-1.251177435e+00 wat=-1.415974246e+00 pat=5.690311985e-6 ute=-0.13298 ua1=6.9609e-10 ub1=-2.456712840e-19 lub1=4.974744624e-25 wub1=6.115299332e-25 pub1=-2.457527824e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos lmin=1.5e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.848188657e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.602615542e-07 wvth0=-4.899759853e-07 pvth0=1.249656648e-12 k1=0.64774 k2=-2.933185363e-01 lk2=3.052625335e-07 wk2=1.021472801e-06 pk2=-1.446301526e-12 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-3.897420539e+05 lvsat=8.053429813e-01 wvsat=3.334604818e+00 pvsat=-5.589086733e-6 ua=-4.785714481e-10 lua=-3.455397567e-15 wua=-1.212718283e-14 pua=1.622766918e-20 ub=-8.352020653e-19 lub=5.423136126e-24 wub=1.840910224e-23 pub=-2.486701119e-29 uc=5.250310988e-11 luc=3.825209488e-17 wuc=-1.773250065e-16 puc=2.044223870e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.219351604e-03 lu0=-1.147085513e-09 wu0=-6.810067359e-09 pu0=4.846124340e-15 a0=-4.931314979e-01 la0=-3.576434503e-07 wa0=1.141731368e-05 pa0=1.067095370e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-8.857177354e-02 lags=1.007675135e-07 wags=1.628309621e-06 pags=3.013259555e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-6.951170377e-03 lpdiblc2=2.875453710e-08 wpdiblc2=2.433040489e-08 ppdiblc2=-5.340206418e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-6.358626674e-03 ldelta=2.194166251e-08 wdelta=1.611990837e-07 pdelta=-6.432210840e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.164150355e-01 lkt1=4.543286592e-07 wkt1=1.561953147e-06 pkt1=-3.153044529e-12 kt2=-2.078416526e-01 lkt2=3.084437267e-07 wkt2=1.060409991e-06 pkt2=-2.140601931e-12 at=-8.494857770e+05 lat=1.641228386e+00 wat=7.328418389e+00 pat=-1.196159993e-5 ute=-0.13298 ua1=8.484518720e-10 lua1=-3.075660548e-16 wua1=-3.238449524e-16 pua1=6.537312324e-22 ub1=3.632596456e-20 lub1=-7.178069341e-26 wub1=-2.446119733e-24 pub1=3.714811963e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos lmin=1e-06 lmax=1.5e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.975234242e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.409677130e-07 wvth0=-2.468313935e-07 pvth0=8.804038984e-13 k1=0.64774 k2=2.810808736e-02 lk2=-1.828736157e-07 wk2=-5.515052775e-07 pk2=9.425094987e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=4.285892796e+05 lvsat=-4.374199901e-01 wvsat=-2.349753621e+00 pvsat=3.043492633e-6 ua=-3.233376441e-09 lua=7.282008095e-16 wua=5.245500136e-16 pua=-2.985948162e-21 ub=3.133821903e-18 lub=-6.044419688e-25 wub=6.855791064e-26 pub=2.985948162e-30 uc=1.043592772e-10 luc=-4.049953287e-17 wuc=-2.431769813e-16 puc=3.044288179e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.754763276e-03 lu0=2.595773874e-09 wu0=2.694701863e-09 pu0=-9.588340963e-15 a0=-2.471102242e+00 la0=2.646211711e-06 wa0=2.292543724e-05 pa0=-1.640977401e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-2.234836086e+00 lags=3.360202543e-06 wags=1.484938024e-05 pags=-1.706498544e-11 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-7.903915549e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.562101358e-07 wvoff=-5.081333947e-07 pvoff=7.716793206e-13 nfactor='2.752212005e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.263771910e-07 wnfactor=-1.061667024e-06 pnfactor=1.612305934e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.736747415e-02 lpdiblc2=-8.177093998e-09 wpdiblc2=-1.180480478e-07 ppdiblc2=1.628216848e-13 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.482887360e-03 ldelta=3.958488016e-09 wdelta=3.045366445e-08 pdelta=1.342350763e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.286908185e-01 lkt1=1.692403384e-07 wkt1=-1.650228519e-07 pkt1=-5.303637942e-13 kt2=5.850083813e-02 lkt2=-9.603862851e-08 wkt2=-1.060409991e-06 pkt2=1.080191940e-12 at=9.476210856e+05 lat=-1.087956936e+00 wat=-5.149513256e+00 pat=6.988073353e-6 ute=3.519795030e-01 lute=-7.364861740e-07 wute=-2.021008904e-06 pute=3.069215277e-12 ua1=5.147883852e-10 lua1=1.991536678e-16 wua1=1.016722379e-15 pua1=-1.382128048e-21 ub1=-9.391785227e-21 lub1=-2.351204106e-27 wub1=-7.648193364e-27 pub1=1.161496709e-32 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos lmin=5e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-7.220578437e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=8.775539610e-08 wvth0=1.127420182e-06 pvth0=-5.194843404e-13 k1=0.64774 k2=-2.197450652e-01 lk2=6.960323742e-08 wk2=7.018996203e-07 pk2=-3.342776675e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-4.290240392e+04 lvsat=4.286737082e-02 wvsat=5.917903168e-01 pvsat=4.707419290e-8 ua=-1.748606390e-09 lua=-7.842676270e-16 wua=-7.200583488e-15 pua=4.883297705e-21 ub=1.449621924e-18 lub=1.111176761e-24 wub=9.495372335e-24 pub=-6.616723486e-30 uc=3.551119815e-11 luc=2.963290707e-17 wuc=2.803981784e-16 puc=-2.289136365e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=5.657598701e-03 lu0=-1.379868946e-09 wu0=-1.563385660e-08 pu0=9.082136754e-15 a0=8.124849089e-01 la0=-6.986307590e-07 wa0=2.546171417e-06 pa0=4.349667016e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.525626381e+00 lags=-4.704113511e-07 wags=-2.453422547e-06 pags=5.606011275e-13 b0=-6.863384714e-07 lb0=6.991421156e-13 wb0=1.434426333e-11 pb0=-1.461185556e-17 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.847608445e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=5.334929131e-08 wvoff=5.081333947e-07 pvoff=-2.635459259e-13 nfactor='2.322387995e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.114651860e-07 wnfactor=1.061667024e-06 pnfactor=-5.506389104e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-4.385445496e-02 lpdiblc2=5.418693020e-08 wpdiblc2=1.335083363e-07 ppdiblc2=-9.342748354e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=4.011694927e-03 ldelta=5.457125545e-09 wdelta=1.165855658e-07 pdelta=4.649638431e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-3.030118372e-01 lkt1=-1.625141843e-07 wkt1=-1.284551785e-06 pkt1=6.100499507e-13 kt2=-1.478799484e-02 lkt2=-2.138259236e-8 at=-3.068657850e+05 lat=1.899323868e-01 wat=3.484991853e+00 pat=-1.807508450e-6 ute=-3.425336980e-01 lute=-2.901682929e-08 wute=2.021008904e-06 pute=-1.048206373e-12 ua1=5.172980422e-10 lua1=1.965971932e-16 wua1=-6.928774262e-16 pua1=3.593643415e-22 ub1=5.977405120e-19 lub1=-6.208095544e-25 wub1=7.648193364e-27 pub1=-3.966773729e-33 uc1=-2.348171346e-11 luc1=1.377294237e-17 puc1=-2.350988702e-38 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos lmin=3.5e-07 lmax=5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.788856617e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.349842807e-08 wvth0=2.037607703e-07 pvth0=-4.042376817e-14 k1=0.64774 k2=-1.031748421e-01 lk2=9.143508357e-09 wk2=1.197847226e-07 pk2=-3.236086522e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=6.861482019e+04 lvsat=-1.497159505e-02 wvsat=1.010442201e+00 pvsat=-1.700617001e-7 ua=-4.186846132e-09 lua=4.803376062e-16 wua=7.657860509e-15 pua=-2.823108566e-21 ub=4.648955398e-18 lub=-5.481735421e-25 wub=-1.127934098e-23 pub=4.158185450e-30 uc=1.651655211e-10 luc=-3.761295578e-17 wuc=-5.565581283e-16 puc=2.051779368e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.581968835e-04 lu0=1.368692304e-09 wu0=1.437906052e-08 pu0=-6.484212771e-15 a0=-4.305909324e+00 la0=1.956050002e-06 wa0=3.780167702e-05 pa0=-1.393577724e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.120307807e+00 lags=-2.601908465e-07 wags=-4.926593924e-06 pags=1.843323828e-12 b0=2.287794905e-06 lb0=-8.434070306e-13 wb0=-4.781421109e-11 pb0=1.762694799e-17 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.723233350e-01 lpdiblc2=1.208179572e-07 wpdiblc2=5.122222396e-07 ppdiblc2=-2.898493431e-13 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=7.317609143e-04 ldelta=7.158279720e-09 wdelta=1.582480458e-07 pdelta=2.488793078e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.025608325e-01 lkt1=-7.151600091e-09 wkt1=-3.745950342e-07 pkt1=1.380963323e-13 kt2=-0.056015 at=1.431951817e+05 lat=-4.349398388e-2 ute=-0.39848 ua1=8.9635e-10 ub1=-5.9922e-19 uc1=3.0734e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.367536275e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=4.996140086e-8 k1=0.64774 k2=-7.405551253e-02 wk2=4.596739352e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.105700400e-09 wua=7.261831520e-16 ub=3.068500280e-18 wub=-5.083282064e-25 uc=3.083053126e-11 wuc=8.849267890e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.283858446e-03 wu0=1.677693674e-9 a0=1.785001752e+00 wa0=-9.520261123e-8 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.807462932e-01 wags=1.241773190e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=7.574465868e-04 wpdiblc2=4.381062956e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.333849813e-02 wdelta=2.154585412e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.60135 kt2=-0.055045 at=2.898042114e+05 wat=-2.076883815e-2 ute=-1.212209238e-01 wute=-5.013568481e-7 ua1=6.8217e-10 ub1=-1.464496940e-19 wub1=-1.082012896e-26 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.367536275e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=4.996140086e-8 k1=0.64774 k2=-7.405551253e-02 wk2=4.596739352e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.105700400e-09 wua=7.261831520e-16 ub=3.068500280e-18 wub=-5.083282064e-25 uc=3.083053126e-11 wuc=8.849267890e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.283858446e-03 wu0=1.677693674e-9 a0=1.785001752e+00 wa0=-9.520261123e-8 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.807462932e-01 wags=1.241773190e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=7.574465868e-04 wpdiblc2=4.381062956e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.333849813e-02 wdelta=2.154585412e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.60135 kt2=-0.055045 at=2.898042114e+05 wat=-2.076883815e-2 ute=-1.212209238e-01 wute=-5.013568481e-7 ua1=6.8217e-10 ub1=-1.464496940e-19 wub1=-1.082012896e-26 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.238555089e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.034255632e-07 wvth0=-3.072902883e-08 pvth0=6.470287175e-13 k1=0.64774 k2=-5.550103971e-02 lk2=-1.487819162e-07 wk2=-5.211272809e-08 pk2=4.547336547e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.150006192e-09 lua=3.552728600e-16 wua=9.450541186e-16 pua=-1.755050771e-21 ub=3.068500280e-18 wub=-5.083282064e-25 uc=3.083053126e-11 wuc=8.849267890e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.968138465e-03 lu0=2.531649603e-09 wu0=3.076738780e-09 pu0=-1.121846003e-14 a0=1.823118512e+00 la0=-3.056451471e-07 wa0=-3.104986854e-07 pa0=1.726384941e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.405866900e-01 lags=3.220260026e-07 wags=-2.727087004e-08 pags=3.182492064e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.486114269e-03 lpdiblc2=1.799034047e-08 wpdiblc2=8.066850034e-09 ppdiblc2=-2.955505498e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.182709075e-02 ldelta=1.211945438e-08 wdelta=5.641230547e-09 pdelta=1.275336893e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.113966375e-01 lkt1=8.056052002e-8 kt2=-0.055045 at=3.076814106e+05 lat=-1.433510927e-01 wat=-4.163453696e-02 pat=1.673148401e-7 ute=-1.094070063e-01 lute=-9.473172904e-08 wute=-1.005051899e-06 pute=4.038956840e-12 ua1=6.681850806e-10 lua1=1.121402439e-16 ub1=-1.711339750e-19 lub1=1.979347329e-25 wub1=-2.169072031e-26 pub1=8.716752161e-32 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.039100293e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.835795644e-07 wvth0=-2.129817265e-08 pvth0=6.091293601e-13 k1=0.64774 k2=-9.931248826e-02 lk2=2.728118053e-08 wk2=9.552123541e-08 pk2=-1.385563109e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.914012137e-09 lua=-5.931058303e-16 wua=7.441788419e-17 pua=1.743735886e-21 ub=2.772825385e-18 lub=1.188215396e-24 wub=3.609583513e-25 pub=-3.493362771e-30 uc=-1.863340926e-12 luc=1.313853929e-16 wuc=2.135424088e-16 puc=-5.025317221e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.353130284e-03 lu0=9.845003037e-10 wu0=9.833575578e-10 pu0=-2.805883116e-15 a0=1.475377148e+00 la0=1.091807427e-06 wa0=1.577245277e-06 pa0=-5.859806772e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.135456361e-02 lags=1.524536684e-06 wags=1.118740464e-06 pags=-4.287174969e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.508014359e-03 lpdiblc2=1.807834938e-08 wpdiblc2=4.344918707e-09 ppdiblc2=-1.459789704e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.265636977e-02 ldelta=8.786868099e-09 wdelta=6.878321653e-09 pdelta=1.225622470e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.59135 kt2=-0.055045 at=2.856943313e+05 lat=-5.499260646e-02 wat=5.445867726e-02 pat=-2.188506357e-7 ute=-0.13298 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos lmin=1.5e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-6.967649991e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.057280846e-07 wvth0=5.570396093e-07 pvth0=-5.583350951e-13 k1=0.64774 k2=-1.022987769e-01 lk2=3.330946704e-08 wk2=7.783366166e-08 pk2=-1.028512017e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=5.227102819e+05 lvsat=-8.053429813e-01 wvsat=-1.172917020e+00 pvsat=2.367714808e-6 ua=-2.999264251e-09 lua=-4.210112242e-16 wua=3.250597813e-16 pua=1.237776367e-21 ub=2.885055096e-18 lub=9.616623286e-25 wub=3.100210220e-26 pub=-2.827294939e-30 uc=-3.421588653e-11 luc=1.966940209e-16 wuc=2.510675296e-16 puc=-5.782819949e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.013714455e-03 lu0=-3.489912352e-10 wu0=-8.542101990e-10 pu0=9.035322237e-16 a0=1.706721084e+00 la0=6.248038337e-07 wa0=5.500243306e-07 pa0=-3.786202072e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.199558772e-01 lags=1.164002249e-06 wags=1.041805580e-07 pags=-2.239128543e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-7.580401644e-03 lpdiblc2=3.033640433e-08 wpdiblc2=2.743881238e-08 ppdiblc2=-6.121650098e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-1.428852753e-02 ldelta=6.317931976e-08 wdelta=2.003728574e-07 pdelta=-2.680364651e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-3.662849645e-01 lkt1=-4.543286592e-07 wkt1=-6.616930048e-07 pkt1=1.335729893e-12 kt2=9.775165259e-02 lkt2=-3.084437267e-07 wkt2=-4.492233810e-07 pkt2=9.068270241e-13 at=1.116542389e+06 lat=-1.732188192e+00 wat=-2.383776478e+00 pat=4.703104952e-6 ute=-0.13298 ua1=9.105019571e-10 lua1=-4.328237693e-16 wua1=-6.303728693e-16 pua1=1.272505344e-21 ub1=-9.541705012e-19 lub1=1.680107382e-24 wub1=2.446940732e-24 pub1=-4.939529143e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos lmin=1e-06 lmax=1.5e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-6.360506158e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.135238827e-07 wvth0=4.374940411e-07 pvth0=-3.767866203e-13 k1=0.64774 k2=-1.320229154e-01 lk2=7.845017851e-08 wk2=2.395431569e-07 pk2=-3.484321352e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-2.981872707e+05 lvsat=4.413171914e-01 wvsat=1.240528351e+00 pvsat=-1.297476073e-6 ua=-3.158226276e-09 lua=-1.796027491e-16 wua=1.533075970e-16 pua=1.498608681e-21 ub=3.626402232e-18 lub=-1.641882068e-25 wub=-2.364792857e-24 pub=8.110910550e-31 uc=1.587879368e-10 luc=-9.641220046e-17 wuc=-5.120549953e-16 puc=5.806378431e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.834873398e-03 lu0=-1.596048370e-09 wu0=-7.581058780e-09 pu0=1.111929446e-14 a0=2.762490622e+00 la0=-9.785458552e-07 wa0=-2.928553380e-06 pa0=1.496557362e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.344193386e+00 lags=-5.433266657e-07 wags=-2.831053988e-06 pags=2.218480077e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='6.811555414e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.491119355e-06 wnfactor=-2.111485594e-05 pnfactor=3.206618154e-11 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.536555663e-02 lpdiblc2=4.215936888e-08 wpdiblc2=4.365338612e-08 ppdiblc2=-8.584084445e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.760430605e-02 ldelta=-1.562799143e-08 wdelta=-1.282264009e-07 pdelta=2.309924415e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.559390125e-01 lkt1=2.892869090e-07 wkt1=9.575850443e-07 pkt1=-1.123394813e-12 kt2=-2.470924670e-01 lkt2=2.152555198e-07 wkt2=4.492233810e-07 pkt2=-4.576036431e-13 at=-6.523731436e+05 lat=9.541842260e-01 wat=2.754471036e+00 pat=-3.100120326e-6 ute=-6.728429516e-01 lute=8.198655707e-07 wute=3.041622220e-06 pute=-4.619174792e-12 ua1=5.929966613e-10 lua1=4.935723577e-17 wua1=6.303728693e-16 pua1=-6.421324751e-22 ub1=4.843913298e-19 lub1=-5.045717358e-25 wub1=-2.446940732e-24 pub1=2.492588411e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos lmin=5e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.729376470e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.263195850e-08 wvth0=-1.032355824e-07 pvth0=1.740303144e-13 k1=0.64774 k2=-2.800167201e-02 lk2=-2.751158113e-08 wk2=-2.453142760e-07 pk2=1.454703131e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=4.449418513e+03 lvsat=1.330348148e-01 wvsat=3.578719351e-01 pvsat=-3.983537016e-7 ua=-3.875550889e-09 lua=5.511035544e-16 wua=3.306539353e-15 pua=-1.713446614e-21 ub=4.018647391e-18 lub=-5.637506993e-25 wub=-3.195634026e-24 pub=1.657431566e-30 uc=7.554278137e-11 luc=-1.161410666e-17 wuc=8.264183708e-17 puc=-2.515305867e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=7.972154451e-04 lu0=1.498277092e-09 wu0=8.376475571e-09 pu0=-5.135927699e-15 a0=1.751874990e+00 la0=5.092281150e-08 wa0=-2.094423101e-06 pa0=6.468663817e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.245152789e+00 lags=-4.424384659e-07 wags=-1.067880759e-06 pags=4.224148505e-13 b0=3.079656446e-06 lb0=-3.137107437e-12 wb0=-4.259781692e-12 pb0=4.339247919e-18 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='4.393102912e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=1.036408595e-5 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.164733796e-02 lpdiblc2=3.837178684e-08 wpdiblc2=-2.559507941e-08 ppdiblc2=-1.530054881e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.407807124e-03 ldelta=2.022509819e-08 wdelta=1.245087844e-07 pdelta=-2.645751870e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.336420617e-01 lkt1=-3.902249140e-08 wkt1=-1.452366304e-07 pkt1=-8.077935669e-28 kt2=-7.101226750e-03 lkt2=-2.921275711e-08 wkt2=-3.797269586e-08 pkt2=3.868107650e-14 at=5.231607620e+05 lat=-2.432792647e-01 wat=-6.153459293e-01 pat=3.325605744e-7 ute=6.276076410e-01 lute=-5.048449276e-07 wute=-2.771497071e-06 pute=1.302388239e-12 ua1=3.770396810e-10 lua1=2.693428935e-16 ub1=5.444703747e-19 lub1=-5.657715553e-25 wub1=2.708030978e-25 pub1=-2.758549296e-31 uc1=-2.348171346e-11 luc1=1.377294237e-17 puc1=-1.175494351e-38 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos lmin=3.5e-07 lmax=5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.513537551e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.196105192e-08 wvth0=6.775293165e-08 pvth0=8.534626665e-14 k1=0.64774 k2=-7.696929515e-02 lk2=-2.114278552e-09 wk2=-9.670888937e-09 pk2=2.325269217e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=5.174240005e+05 lvsat=-1.330220170e-01 wvsat=-1.206678740e+00 pvsat=4.131083288e-7 ua=-2.884741227e-09 lua=3.721516887e-17 wua=1.225451860e-15 pua=-6.340801806e-22 ub=2.706020166e-18 lub=1.170499744e-25 wub=-1.681225393e-24 pub=8.719759564e-31 uc=-1.699849067e-11 luc=3.638288679e-17 wuc=3.433335470e-16 puc=-1.603621175e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.909127265e-03 lu0=-1.157315329e-10 wu0=-3.162563975e-09 pu0=8.488528573e-16 a0=5.723981007e+00 la0=-2.009229834e-06 wa0=-1.174606145e-05 pa0=5.652736872e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-1.458064201e-01 lags=2.789894827e-07 wags=1.328020489e-06 pags=-8.202313110e-13 b0=-1.026552149e-05 lb0=3.784435823e-12 wb0=1.419927231e-11 pb0=-5.234632732e-18 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='4.393102912e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=1.036408595e-5 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-3.803039963e-02 lpdiblc2=5.205549369e-08 wpdiblc2=-1.511859353e-07 ppdiblc2=4.983777653e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=6.008926949e-02 ldelta=-9.691680674e-09 wdelta=-1.349785214e-07 pdelta=1.081268699e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.851178723e-01 lkt1=3.954119515e-08 wkt1=3.323740287e-08 pkt1=-9.256644972e-14 kt2=-8.163756030e-02 lkt2=9.445884967e-09 wkt2=1.265756529e-07 pkt2=-4.666274731e-14 at=1.251002968e+05 lat=-3.682321410e-02 wat=8.938887605e-02 pat=-3.295365610e-8 ute=-2.162096147e-01 lute=-6.719488890e-08 wute=-9.004171616e-07 pute=3.319432887e-13 ua1=8.9635e-10 ub1=-4.164921597e-19 lub1=-6.736353195e-26 wub1=-9.026769927e-25 pub1=3.327763868e-31 uc1=3.0734e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.391420250e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=5.698330842e-8 k1=0.64774 k2=-7.427707519e-02 wk2=5.248135345e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.845727890e-09 wua=-3.813810835e-17 ub=2.874731822e-18 wub=6.135260909e-26 uc=5.921166538e-11 wuc=5.051917541e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.058205904e-03 wu0=-5.988940464e-10 a0=1.905731793e+00 wa0=-4.501498965e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.696666698e-01 wags=4.499191333e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.649641422e-03 wpdiblc2=-1.182004996e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.431423104e-02 wdelta=-1.072288844e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.919499200e-01 wkt1=-2.763631040e-8 kt2=-0.055045 at=2.867256339e+05 wat=-1.171779561e-2 ute=-0.29175 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.391420250e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=5.698330842e-8 k1=0.64774 k2=-7.427707519e-02 wk2=5.248135345e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.845727890e-09 wua=-3.813810835e-17 ub=2.874731822e-18 wub=6.135260909e-26 uc=5.921166538e-11 wuc=5.051917541e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.058205904e-03 wu0=-5.988940464e-10 a0=1.905731793e+00 wa0=-4.501498965e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.696666698e-01 wags=4.499191333e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.649641422e-03 wpdiblc2=-1.182004996e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.431423104e-02 wdelta=-1.072288844e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.919499200e-01 wkt1=-2.763631040e-8 kt2=-0.055045 at=2.867256339e+05 wat=-1.171779561e-2 ute=-0.29175 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.505853397e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=9.175999280e-08 wvth0=4.785688742e-08 pvth0=7.318162131e-14 k1=0.64774 k2=-7.232563365e-02 lk2=-1.564793646e-08 wk2=-2.648287320e-09 pk2=6.331868908e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.825031897e-09 lua=-1.659540268e-16 wua=-1.037290911e-17 pua=-2.226395537e-22 ub=2.913924089e-18 lub=-3.142692632e-25 wub=-5.387296777e-26 pub=9.239541480e-31 uc=5.921166538e-11 wuc=5.051917541e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.291267286e-03 lu0=-1.868838816e-09 wu0=-8.132705380e-10 pu0=1.719011126e-15 a0=1.905230760e+00 la0=4.017607915e-09 wa0=-5.519093517e-07 pa0=8.159739644e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.013789474e-01 lags=5.475756865e-07 wags=8.800020696e-08 pags=-3.448686687e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.699474560e-03 lpdiblc2=-3.995947414e-10 wpdiblc2=-4.238814607e-09 ppdiblc2=2.451150167e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.874169419e-02 ldelta=4.468425049e-08 wdelta=-1.468775889e-08 pdelta=3.179292827e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.925526379e-01 lkt1=4.832986717e-09 wkt1=-5.540150964e-08 pkt1=2.226395537e-13 kt2=-0.055045 at=3.015098979e+05 lat=-1.185499121e-01 wat=-2.349024009e-02 pat=9.439917078e-8 ute=-4.512604636e-01 lute=1.279059376e-6 ua1=6.681850806e-10 lua1=1.121402439e-16 ub1=-1.549156456e-19 lub1=3.837444072e-26 wub1=-6.937273857e-26 pub1=5.562760570e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.366569820e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.578672855e-08 wvth0=7.497813008e-08 pvth0=-3.580929610e-14 k1=0.64774 k2=-7.158490117e-02 lk2=-1.862468475e-08 wk2=1.400190755e-08 pk2=-3.592699766e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.842608411e-09 lua=-9.532007783e-17 wua=-1.355096390e-16 pua=2.802417914e-22 ub=2.807021019e-18 lub=1.153372942e-25 wub=2.604229137e-25 pub=-3.390925676e-31 uc=7.367640742e-11 luc=-5.812880793e-17 wuc=-8.545055696e-18 puc=5.464154449e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.865507701e-03 lu0=-1.578579308e-10 wu0=-5.230361450e-10 pu0=5.526592320e-16 a0=2.194314136e+00 la0=-1.157708743e-06 wa0=-5.364352195e-07 pa0=7.537887657e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.052144290e-01 lags=1.302967090e-07 wags=4.898954833e-08 pags=-1.880982904e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-2.425186950e-05 lpdiblc2=1.054612209e-08 wpdiblc2=-1.735488266e-11 ppdiblc2=7.546911442e-15 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.206358510e-02 ldelta=7.152126696e-08 wdelta=8.621113313e-09 pdelta=-6.187738754e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.59135 kt2=-0.055045 at=3.042176405e+05 lat=-1.294313956e-1 ute=-1.430749758e-01 lute=4.056822513e-08 wute=2.967930972e-08 pute=-1.192709064e-13 ua1=6.9609e-10 ub1=-1.690722107e-19 lub1=9.526479219e-26 wub1=1.387454771e-25 pub1=-2.800792512e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos lmin=1.5e-06 lmax=2e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.304483089e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.325355966e-08 wvth0=6.806720970e-08 pvth0=-2.185853211e-14 k1=0.64774 k2=-7.959227919e-02 lk2=-2.460551081e-09 wk2=1.107637670e-08 pk2=2.312937700e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.889828010e-09 wua=3.316357248e-18 ub=2.864156732e-18 wub=9.244345829e-26 uc=4.488059638e-11 wuc=1.852323705e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.817651315e-03 lu0=-6.125239980e-11 wu0=-2.777830006e-10 pu0=5.757774583e-17 a0=2.103624126e+00 la0=-9.746369013e-07 wa0=-6.168737881e-07 pa0=9.161664843e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.767321073e-01 lags=5.915236902e-07 wags=2.312587873e-07 pags=-5.560370010e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.728487182e-03 lpdiblc2=1.398638523e-08 wpdiblc2=1.023413705e-08 ppdiblc2=-1.314731400e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=6.787581986e-02 ldelta=-4.114437979e-08 wdelta=-4.119098122e-08 pdelta=3.867604616e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.59135 kt2=-0.055045 at=3.365855781e+05 lat=-1.947710947e-01 wat=-9.069721532e-02 pat=1.830863872e-7 ute=-1.229783149e-01 wute=-2.940503427e-8 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos lmin=1e-06 lmax=1.5e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.898660706e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.837685944e-08 wvth0=7.710309000e-09 pvth0=6.980277692e-14 k1=0.64774 k2=-4.724474936e-02 lk2=-5.158528898e-08 wk2=-9.705329339e-09 pk2=3.387317949e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.209378915e-09 lua=4.852875807e-16 wua=3.036967650e-16 pua=-4.561742082e-22 ub=2.756042508e-18 lub=1.641882068e-25 wub=1.940716937e-25 pub=-1.543382279e-31 uc=-5.296427373e-11 luc=1.485926012e-16 wuc=1.104981977e-16 puc=-1.396782339e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=7.072912728e-04 lu0=3.143656431e-09 wu0=1.614057688e-09 pu0=-2.815475576e-15 a0=1.812442528e+00 la0=-5.324325126e-07 wa0=-1.354043833e-07 pa0=1.849805653e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.574549773e-01 lags=1.652025000e-07 wags=-2.240359718e-07 pags=1.353986614e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='-1.736955414e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=6.491119355e-06 wnfactor=4.017834283e-06 pnfactor=-6.101704123e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=3.178277226e-03 lpdiblc2=6.534702924e-09 wpdiblc2=-1.086563376e-08 ppdiblc2=1.889595844e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.596066583e-03 ldelta=5.951169892e-08 wdelta=-2.236188875e-08 pdelta=1.008115073e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.263239211e-01 lkt1=-9.875217986e-08 wkt1=-1.148596123e-08 pkt1=1.744321246e-14 kt2=-9.429581446e-02 lkt2=5.960844563e-08 wkt2=-2.646977960e-23 at=2.329199329e+05 lat=-3.733874421e-02 wat=1.517023084e-01 pat=-1.850348616e-7 ute=5.998369705e-01 lute=-1.097707047e-06 wute=-7.000669325e-07 pute=1.018504045e-12 ua1=8.074086184e-10 lua1=-1.690545764e-16 ub1=-3.478991714e-19 lub1=3.432451447e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos lmin=5e-07 lmax=1e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.530446239e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.598028971e-08 wvth0=1.322795706e-07 pvth0=-5.709032423e-14 k1=0.64774 k2=-1.292466637e-01 lk2=3.194637108e-08 wk2=5.234680956e-08 pk2=-2.933654206e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.191582443e+05 lvsat=4.687601412e-03 wvsat=2.062706953e-02 pvsat=-2.101186752e-8 ua=-2.706734681e-09 lua=-2.673348149e-17 wua=-1.297896482e-16 pua=-1.460110594e-23 ub=2.956227065e-18 lub=-3.973079241e-26 wub=-7.210976655e-26 pub=1.168088475e-31 uc=1.182349972e-10 luc=-2.580039207e-17 wuc=-4.287361885e-17 puc=1.655473392e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.189104848e-03 lu0=-4.031103765e-10 wu0=-1.595706408e-09 pu0=4.541666703e-16 a0=8.128616885e-01 la0=4.857955078e-07 wa0=6.662835187e-07 pa0=-6.316628245e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=9.212092706e-01 lags=-3.072031296e-07 wags=-1.154842234e-07 pags=2.482188010e-14 b0=2.235533608e-06 lb0=-2.277237487e-12 wb0=-1.778053795e-12 pb0=1.811223389e-18 b1=1.018421991e-07 lb1=-1.037420653e-13 wb1=-2.994168801e-13 pb1=3.050025020e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='4.635289709e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=-1.972127110e-6 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-2.277765037e-02 lpdiblc2=3.297483835e-08 wpdiblc2=7.128128137e-09 ppdiblc2=5.665229105e-16 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.116756451e-02 ldelta=9.015444693e-09 wdelta=-1.884529238e-08 pdelta=6.498952255e-15 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.771981236e-01 lkt1=-4.692891909e-08 wkt1=-1.718145991e-08 pkt1=2.324496066e-14 kt2=-2.001707455e-02 lkt2=-1.605596417e-8 at=3.335427455e+05 lat=-1.398386754e-01 wat=-5.786744388e-02 pat=2.844441448e-8 ute=-4.254045488e-01 lute=-5.333964737e-08 wute=3.243671907e-07 pute=-2.504089669e-14 ua1=3.770396810e-10 lua1=2.693428935e-16 ub1=6.365800213e-19 lub1=-6.595995073e-25 wub1=3.443831106e-41 pub1=3.831675488e-47 uc1=-2.348171346e-11 luc1=1.377294237e-17 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos lmin=3.5e-07 lmax=5e-07 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.721210613e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.587437935e-08 wvth0=1.288089778e-07 pvth0=-5.529028396e-14 k1=0.64774 k2=-8.395695939e-02 lk2=8.456639483e-09 wk2=1.087289985e-08 pk2=-7.825891418e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.098155150e+05 lvsat=9.533254674e-03 wvsat=-8.306531983e-03 pvsat=-6.005310421e-9 ua=-2.298687660e-09 lua=-2.383691095e-16 wua=-4.975503143e-16 pua=1.761398023e-22 ub=1.964392279e-18 lub=4.746892784e-25 wub=4.991665272e-25 pub=-1.794864586e-31 uc=1.199657769e-10 luc=-2.669806963e-17 wuc=-5.934249532e-17 puc=2.509639904e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.110444347e-03 lu0=1.563422855e-10 wu0=-8.144298070e-10 pu0=4.895365457e-17 a0=1.994770598e+00 la0=-1.272074574e-07 wa0=-7.821530183e-07 pa0=1.195760276e-13 keta=-1.170787773e-02 lketa=-4.523305745e-10 wketa=-2.564046443e-09 pketa=1.329855508e-15 a1=0.0 a2=0.46703705 ags=3.289019958e-01 wags=-6.762605155e-8 b0=-7.923591064e-06 lb0=2.991843319e-12 wb0=7.313978129e-12 pb0=-2.904404429e-18 b1=-1.058029858e-07 lb1=3.954148069e-15 wb1=3.110616248e-13 pb1=-1.162522696e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='4.635289709e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=-1.972127110e-6 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.055652710e-01 lpdiblc2=7.591305174e-08 wpdiblc2=4.736712695e-08 ppdiblc2=-2.030363502e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-1.964677107e-02 ldelta=4.574365391e-08 wdelta=9.944607568e-08 pdelta=-5.485345725e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.781301771e-01 lkt1=5.419995134e-09 wkt1=1.269352318e-08 pkt1=7.750151303e-15 kt2=-7.245773213e-02 lkt2=1.114264509e-08 wkt2=9.958688462e-08 pkt2=-5.165123564e-14 at=1.571456507e+05 lat=-4.834944024e-02 wat=-4.824720815e-03 pat=9.335409525e-10 ute=-6.321705323e-01 lute=5.390056380e-08 wute=3.225112639e-07 pute=-2.407831098e-14 ua1=6.963047891e-10 lua1=1.037544489e-16 wua1=5.881345205e-16 pua1=-3.050389097e-22 ub1=-2.998808163e-19 lub1=-1.738994116e-25 wub1=-1.245515275e-24 pub1=6.459927251e-31 uc1=3.417709198e-11 luc1=-1.613208536e-17 wuc1=-9.144510324e-17 puc1=4.742846002e-23 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.168079584e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=3.598910718e-8 k1=0.64774 k2=-8.905546576e-02 wk2=1.913994071e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.729170768e-09 wua=-1.477027351e-16 ub=2.790819787e-18 wub=1.402305940e-25 uc=6.950894704e-11 wuc=-4.627609601e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.560156448e-03 wu0=-1.307235739e-10 a0=1.103396541e+00 wa0=3.040516587e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.840456075e-01 wags=-1.565260031e-7 b0=1.932591552e-07 wb0=-1.816651520e-13 b1=-2.220062912e-07 wb1=2.086876898e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.436766387e-03 wpdiblc2=-9.819007605e-10 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.218069925e-02 wdelta=6.827285123e-10 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.634201653e-01 wkt1=-5.445450803e-8 kt2=-0.055045 at=2.656031920e+05 wat=8.137468774e-3 ute=-2.980983259e-01 wute=5.967477101e-9 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos lmin=8e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.168079584e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=3.598910718e-8 k1=0.64774 k2=-8.905546576e-02 wk2=1.913994071e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.729170768e-09 wua=-1.477027351e-16 ub=2.790819787e-18 wub=1.402305940e-25 uc=6.950894704e-11 wuc=-4.627609601e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.560156448e-03 wu0=-1.307235739e-10 a0=1.103396541e+00 wa0=3.040516587e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.840456075e-01 wags=-1.565260031e-7 b0=1.932591552e-07 wb0=-1.816651520e-13 b1=-2.220062912e-07 wb1=2.086876898e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.436766387e-03 wpdiblc2=-9.819007605e-10 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.218069925e-02 wdelta=6.827285123e-10 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.634201653e-01 wkt1=-5.445450803e-8 kt2=-0.055045 at=2.656031920e+05 wat=8.137468774e-3 ute=-2.980983259e-01 wute=5.967477101e-9 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos lmin=4e-06 lmax=8e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.640320008e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=3.786733039e-07 wvth0=6.049685648e-08 pvth0=-1.965191865e-13 k1=0.64774 k2=-1.087788170e-01 lk2=1.581547493e-07 wk2=3.161799668e-08 pk2=-1.000572259e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.668325925e-09 lua=-4.878938008e-16 wua=-1.576777757e-16 pua=7.998640939e-23 ub=2.650326676e-18 lub=1.126565788e-24 wub=1.939107095e-25 pub=-4.304423268e-31 uc=6.359486383e-11 luc=4.742299289e-17 wuc=9.316759271e-19 puc=-4.457799270e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.391716001e-03 lu0=1.350665834e-09 wu0=3.231486594e-11 pu0=-1.307349000e-15 a0=8.384753238e-01 la0=2.124311846e-06 wa0=4.508492927e-07 pa0=-1.177119581e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.080260702e-01 lags=6.095744425e-07 wags=-1.062497417e-07 pags=-4.031479954e-13 b0=-2.227778036e-08 lb0=1.728316326e-12 wb0=2.094129176e-14 pb0=-1.624631173e-18 b1=-2.270386225e-07 lb1=4.035252817e-14 wb1=2.134181214e-13 pb1=-3.793169930e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.359353681e-03 lpdiblc2=3.043977717e-08 wpdiblc2=-4.234835893e-10 ppdiblc2=-4.477754642e-15 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-3.370674291e-03 ldelta=1.247010992e-07 wdelta=6.098044382e-09 pdelta=-4.342354968e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.935819575e-01 lkt1=2.418570058e-07 wkt1=-5.443394093e-08 pkt1=-1.649204317e-16 kt2=-0.055045 at=2.561580453e+05 lat=7.573737243e-02 wat=1.914086410e-02 pat=-8.823243098e-8 ute=-4.232532828e-01 lute=1.003574421e-06 wute=-2.632697401e-08 pute=2.589580619e-13 ua1=6.681850806e-10 lua1=1.121402439e-16 ub1=-2.833833304e-19 lub1=1.068512484e-24 wub1=5.138791290e-26 pub1=-4.120619447e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos lmin=2e-06 lmax=4e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.505106779e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-7.752972820e-08 wvth0=-6.000084965e-09 pvth0=7.070907978e-14 k1=0.64774 k2=-5.383108123e-02 lk2=-6.266124394e-08 wk2=-2.686825230e-09 pk2=3.780201817e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.906143344e-09 lua=4.678123584e-16 wua=-7.578629386e-17 pua=-2.491072037e-22 ub=3.080199636e-18 lub=-6.009453324e-25 wub=3.632828354e-27 pub=3.342188317e-31 uc=7.539557648e-11 wuc=-1.016108837e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.545867443e-03 lu0=7.311843720e-10 wu0=-2.225717455e-10 pu0=-2.830476451e-16 a0=1.552040238e+00 la0=-7.432593660e-07 wa0=6.730738206e-08 pa0=3.642030354e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=7.849888296e-01 lags=-5.034433352e-07 wags=-3.080014264e-07 pags=4.076224210e-13 b0=5.928558493e-07 lb0=-7.436935105e-13 wb0=-5.572892412e-13 pb0=6.990778494e-19 b1=-2.143595683e-07 lb1=-1.060021633e-14 wb1=2.014997090e-13 pb1=9.964288149e-21 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.049443446e-03 lpdiblc2=2.075965255e-08 wpdiblc2=-1.026637069e-09 ppdiblc2=-2.053888895e-15 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.184251420e-02 ldelta=-1.680855675e-08 wdelta=-9.971238266e-09 pdelta=2.115335338e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.333983872e-01 wkt1=-5.447497964e-8 kt2=-0.055045 at=3.014640320e+05 lat=-1.063317576e-01 wat=2.588413997e-03 pat=-2.171384459e-8 ute=-1.286577915e-01 lute=-1.803032228e-07 wute=1.612704115e-08 pute=8.835002159e-14 ua1=6.9609e-10 ub1=8.786315888e-20 lub1=-4.233990764e-25 wub1=-1.027758258e-25 pub1=2.074689346e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos lmin=1.5e-06 lmax=2e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.889173042e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=2.902773295e-8 k1=0.64774 k2=-8.487216747e-02 wk2=1.603951392e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.674398763e-09 wua=-1.991888583e-16 ub=2.782503728e-18 wub=1.691979357e-25 uc=7.539557648e-11 wuc=-1.016108837e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.908081081e-03 wu0=-3.627877036e-10 a0=1.183844897e+00 wa0=2.477260447e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.355933979e-01 wags=-1.060736967e-7 b0=2.244454421e-07 wb0=-2.109805112e-13 b1=-2.196106965e-07 wb1=2.064358116e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.133334661e-02 wpdiblc2=-2.044091213e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.351590229e-02 wdelta=5.076961650e-10 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.333983872e-01 wkt1=-5.447497964e-8 kt2=-0.055045 at=2.487894752e+05 wat=-8.168176204e-3 ute=-2.179762847e-01 wute=5.989381734e-8 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos lmin=1e-06 lmax=1.5e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.855062759e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=1.466853249e-07 wvth0=9.761286706e-08 pvth0=-1.041571568e-13 k1=0.64774 k2=-1.149461471e-01 lk2=4.567199954e-08 wk2=5.393452615e-08 pk2=-5.754944979e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=5.656787592e+04 lvsat=1.020416552e-01 wvsat=6.316113417e-02 pvsat=-9.591997221e-8 ua=-1.980692437e-09 lua=-1.053500580e-15 wua=-8.512783543e-16 pua=9.902989736e-22 ub=2.035998520e-18 lub=1.133683867e-24 wub=8.709188036e-25 pub=-1.065671905e-30 uc=1.161816040e-10 luc=-6.193990461e-17 wuc=-4.850028051e-17 puc=5.822400585e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.190995380e-03 lu0=-1.948304215e-09 wu0=-1.660652042e-09 pu0=1.971008167e-15 a0=8.227061687e-01 la0=5.484451361e-07 wa0=7.949557127e-07 pa0=-8.310530715e-13 keta=-1.090507747e-02 lketa=-2.543629479e-09 wketa=-1.574440580e-09 pketa=2.391032060e-15 a1=0.0 a2=0.46703705 ags=4.449494350e-01 lags=1.376569074e-07 wags=-2.122806620e-07 pags=1.612917388e-13 b0=3.121958538e-07 lb0=-1.332626014e-13 wb0=-2.934666001e-13 pb0=1.252679114e-19 b1=3.465574884e-07 lb1=-8.598141449e-13 wb1=-3.257668116e-13 pb1=8.082321748e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=3.594807230e-03 lpdiblc2=1.175217153e-08 wpdiblc2=-1.125717530e-08 ppdiblc2=1.399149621e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-5.797965374e-02 ldelta=1.237636337e-07 wdelta=3.363976496e-08 pdelta=-5.031618194e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-2.758292593e-01 lkt1=-3.911586439e-07 wkt1=-2.469529473e-07 pkt1=2.923076280e-13 kt2=-2.042417227e-01 lkt2=2.265783489e-07 wkt2=1.033500333e-07 pkt2=-1.569530449e-13 at=3.013888969e+05 lat=-7.988037476e-02 wat=8.734093450e-02 pat=-1.450453885e-7 ute=-2.078796358e-01 lute=-1.533332632e-08 wute=5.919313915e-08 pute=1.064088440e-15 ua1=9.886995712e-10 lua1=-4.443729884e-16 wua1=-1.704149460e-16 pua1=2.588015098e-22 ub1=-5.320474755e-19 lub1=6.229028876e-25 wub1=1.731008791e-25 pub1=-2.628805155e-31 uc1=7.869009847e-11 luc1=-1.346304339e-16 wuc1=-8.333274177e-17 puc1=1.265536849e-22 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos lmin=5e-07 lmax=1e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.260387295e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.575708859e-08 wvth0=1.289301382e-08 pvth0=-1.785685473e-14 k1=0.64774 k2=-6.635938509e-02 lk2=-3.821148519e-09 wk2=-6.767735454e-09 pk2=4.285212504e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.827200985e+05 lvsat=-2.646393707e-02 wvsat=-3.912158185e-02 pvsat=8.270827870e-9 ua=-3.083649974e-09 lua=7.003262943e-17 wua=2.245137420e-16 pua=-1.055620243e-22 ub=3.301104953e-18 lub=-1.550231268e-25 wub=-3.962977407e-25 pub=2.251845642e-31 uc=6.605715941e-11 luc=-1.088038852e-17 wuc=6.173966047e-18 puc=2.529811218e-24 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.289055168e-03 lu0=-1.088330837e-11 wu0=1.903554908e-10 pu0=8.547008842e-17 a0=1.566917440e+00 la0=-2.096493962e-07 wa0=-4.253491989e-08 pa0=2.206094888e-14 keta=-1.340212453e-02 wketa=7.728036383e-10 a1=0.0 a2=0.46703705 ags=1.189788459e+00 lags=-6.210770888e-07 wags=-3.679508093e-07 pags=3.198659127e-13 b0=5.933804351e-07 lb0=-4.196926811e-13 wb0=-2.344166757e-13 pb0=6.511641061e-20 b1=-9.199840112e-07 lb1=4.303546864e-13 wb1=6.611079322e-13 pb1=-1.970527174e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.054530457e-02 lpdiblc2=4.672012659e-09 wpdiblc2=-2.419571609e-08 ppdiblc2=2.717140549e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.437755642e-02 ldelta=2.968349973e-08 wdelta=-3.062550458e-09 pdelta=-1.292918482e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.527032332e-01 lkt1=-7.254086091e-09 wkt1=5.379394710e-08 pkt1=-1.404969976e-14 kt2=5.111240555e-02 lkt2=-3.353941059e-08 wkt2=-6.686228033e-08 pkt2=1.643457951e-14 at=4.359437446e+05 lat=-2.169453431e-01 wat=-1.541252022e-01 pat=1.009252989e-7 ute=-5.892375205e-02 lute=-1.670679821e-07 wute=-2.012769011e-08 pute=8.186464777e-14 ua1=1.360691054e-13 lua1=5.626321659e-16 wua1=3.542924104e-16 pua1=-2.756942623e-22 ub1=1.223079551e-18 lub1=-1.164966034e-24 wub1=-5.513142501e-25 pub1=4.750485779e-31 uc1=-8.171830780e-11 luc1=2.877039114e-17 wuc1=5.474286457e-17 puc1=-1.409772182e-23 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos lmin=3.5e-07 lmax=5e-07 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.194136917e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.229241976e-07 wvth0=-2.027387712e-07 pvth0=9.398164874e-14 k1=0.64774 k2=-2.760129833e-02 lk2=-2.392322400e-08 wk2=-4.210187239e-08 pk2=2.261143930e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=2.180127419e+05 lvsat=-4.476864305e-02 wvsat=-1.100127908e-01 pvsat=4.503890786e-8 ua=-3.063875819e-09 lua=5.977666504e-17 wua=2.217326766e-16 pua=-1.041196108e-22 ub=2.578231905e-18 lub=2.198985938e-25 wub=-7.784763241e-26 pub=6.001882330e-32 uc=1.770416442e-11 luc=1.419813410e-17 wuc=3.678423850e-17 puc=-1.334635964e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.816741375e-04 lu0=9.265239002e-10 wu0=1.656635220e-09 pu0=-6.750232247e-16 a0=1.1627 keta=-1.727822350e-02 lketa=2.010358109e-09 wketa=2.672123140e-09 pketa=-9.850915563e-16 a1=0.0 a2=0.46703705 ags=-7.062579062e-01 lags=3.623168389e-07 wags=9.054325375e-07 pags=-3.405807271e-13 b0=1.350724194e-06 lb0=-8.124928084e-13 wb0=-1.403952408e-12 pb0=6.717019657e-19 b1=-1.350535301e-06 lb1=6.536622654e-13 wb1=1.481119959e-12 pb1=-6.223560549e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-8.378519310e-03 lpdiblc2=1.448694853e-08 wpdiblc2=-4.398919716e-08 ppdiblc2=3.743739341e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.491858311e-01 ldelta=-2.986238598e-08 wdelta=-5.925792104e-08 pdelta=1.621682510e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.896203904e-01 lkt1=6.375868209e-08 wkt1=1.174952156e-07 pkt1=-4.708868115e-14 kt2=1.628729544e-01 lkt2=-9.150457803e-08 wkt2=-1.216258433e-07 pkt2=4.483797527e-14 at=-3.155427851e+04 lat=2.552484406e-02 wat=1.725547223e-01 pat=-6.850887728e-8 ute=-7.956346097e-01 lute=2.150307878e-07 wute=4.761688044e-07 pute=-1.755420106e-13 ua1=1.974016683e-09 lua1=-4.611308839e-16 wua1=-6.129248814e-16 pua1=2.259578221e-22 ub1=-2.966056543e-18 lub1=1.007750347e-24 wub1=1.260711237e-24 pub1=-4.647675010e-31 uc1=-1.644857853e-10 luc1=7.169815716e-17 wuc1=9.529959066e-17 puc1=-3.513267059e-23 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.958567050e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=2.572282540e-8 k1=0.64774 k2=-6.193064985e-02 wk2=5.848563910e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.318606400e-09 wua=1.411254401e-16 ub=3.612858062e-18 wub=-2.625747370e-25 uc=5.989884246e-11 wuc=8.141852311e-20 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.328847096e-03 wu0=-1.738014073e-11 a0=2.006644745e+00 wa0=-1.385471868e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.752969040e-01 wags=-1.522390685e-7 b0=-2.984149951e-07 wb0=5.925911507e-14 b1=2.037138425e-07 wb1=8.141852311e-17 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-3.987916076e-01 wpclm=2.101588488e-7 pdiblc1=0.0 pdiblc2=1.263679999e-03 wpdiblc2=-4.070790458e-10 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.067732025e-02 wdelta=1.419396253e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.407075385e-01 wkt1=8.141852311e-8 kt2=-0.055045 at=2.601941262e+05 wat=1.078795431e-2 ute=-5.868036092e-01 wute=1.474353756e-7 ua1=6.8217e-10 ub1=-7.945766031e-20 wub1=-3.463001183e-26 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.467972681e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=1.019761558e-06 wvth0=5.068410885e-08 pvth0=-4.996913217e-13 k1=0.64774 k2=-8.038753652e-02 lk2=3.694820467e-07 wk2=1.489258604e-08 pk2=-1.810491588e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.318606400e-09 wua=1.411254401e-16 ub=3.612858062e-18 wub=-2.625747370e-25 uc=5.989884246e-11 wuc=8.141852311e-20 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.522592592e-03 lu0=-3.878524244e-09 wu0=-1.123169838e-10 pu0=1.900507908e-15 a0=1.694095300e+00 la0=6.256819500e-06 wa0=1.460454138e-08 pa0=-3.065891610e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.752969040e-01 wags=-1.522390685e-7 b0=-2.525781109e-07 lb0=-9.175927710e-13 wb0=3.679867512e-14 pb0=4.496277985e-19 b1=1.996797525e-07 lb1=8.075705453e-14 wb1=2.058154861e-15 pb1=-3.957160278e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-3.987916076e-01 wpclm=2.101588488e-7 pdiblc1=0.0 pdiblc2=3.280854499e-03 lpdiblc2=-4.038112038e-08 wpdiblc2=-1.395510688e-09 ppdiblc2=1.978707204e-14 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.100496056e-02 ldelta=-2.067454685e-07 wdelta=-3.641230124e-09 pdelta=1.013069335e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.407075385e-01 wkt1=8.141852311e-8 kt2=-0.055045 at=2.298089167e+05 lat=6.082710254e-01 wat=2.567695003e-02 pat=-2.980576686e-7 ute=-5.868036092e-01 wute=1.474353756e-7 ua1=6.8217e-10 ub1=-3.223290114e-20 lub1=-9.453761613e-25 wub1=-5.777052162e-26 pub1=4.632418820e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.042793498e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.230404600e-07 wvth0=-1.778322055e-08 pvth0=4.932457158e-14 k1=0.64774 k2=-1.555012570e-02 lk2=-1.504267817e-07 wk2=-1.406480790e-08 pk2=5.115019291e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.360750016e-09 lua=3.379351207e-16 wua=1.816155682e-16 pua=-3.246763688e-22 ub=3.917726875e-18 lub=-2.444637833e-24 wub=-4.271255273e-25 pub=1.319476017e-30 uc=9.710008322e-11 luc=-2.983039152e-16 wuc=-1.548614961e-17 puc=1.248309581e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.977837869e-03 lu0=-7.528979064e-09 wu0=-2.548895385e-10 pu0=3.043748036e-15 a0=2.793102510e+00 la0=-2.555740160e-06 wa0=-5.069336656e-07 pa0=1.116143342e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=6.754975198e-01 lags=-8.034741687e-07 wags=-1.883120917e-07 pags=2.892571285e-13 b0=2.490386438e-07 lb0=-4.939884469e-12 wb0=-1.120059266e-13 pb0=1.642840562e-18 b1=2.360735722e-07 lb1=-2.110724294e-13 wb1=-1.351055885e-14 pb1=8.526854129e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-3.987916076e-01 wpclm=2.101588488e-7 pdiblc1=0.0 pdiblc2=1.161819637e-03 lpdiblc2=-2.338931089e-08 wpdiblc2=-1.658878685e-09 ppdiblc2=2.189892914e-14 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-2.631295116e-03 ldelta=-1.721448871e-08 wdelta=5.735742671e-09 pdelta=2.611622374e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-9.542935855e-01 lkt1=9.108073242e-07 wkt1=1.223176425e-07 pkt1=-3.279559280e-13 kt2=-0.055045 at=3.422415997e+05 lat=-2.932878707e-01 wat=-2.304076621e-02 pat=9.259289035e-8 ute=-1.080151388e+00 lute=3.955985636e-06 wute=2.955583529e-07 pute=-1.187747053e-12 ua1=6.681850806e-10 lua1=1.121402439e-16 ub1=-1.785117509e-19 lub1=2.275834691e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-4.926732021e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=2.321839366e-07 wvth0=1.465988921e-08 pvth0=-8.105309368e-14 k1=0.64774 k2=-6.544989024e-02 lk2=5.010315652e-08 wk2=3.006484135e-09 pk2=-1.745344018e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.238613915e-09 lua=-1.528877355e-16 wua=8.712694538e-17 pua=5.504080788e-23 ub=3.233315472e-18 lub=3.057754710e-25 wub=-7.139515658e-26 pub=-1.100816158e-31 uc=2.287029360e-11 wuc=1.557672045e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=7.750017662e-04 lu0=1.323459257e-09 wu0=6.451666030e-10 pu0=-5.732670767e-16 a0=1.968183164e+00 la0=7.593260952e-07 wa0=-1.366059806e-07 pa0=-3.720758612e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.208834747e-01 lags=6.215973368e-07 wags=-8.058608961e-08 pags=-1.436565086e-13 b0=-1.645166440e-06 lb0=2.672272263e-12 wb0=5.393595849e-13 pb0=-9.747727075e-19 b1=2.457233235e-07 lb1=-2.498514507e-13 wb1=-2.394458857e-14 pb1=1.271993070e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-3.987916076e-01 wpclm=2.101588488e-7 pdiblc1=0.0 pdiblc2=-1.527591177e-02 lpdiblc2=4.266826062e-08 wpdiblc2=6.972917590e-09 ppdiblc2=-1.278928212e-14 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-4.223357820e-02 ldelta=1.419334242e-07 wdelta=2.632663962e-08 pdelta=-5.663148722e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.869238288e-01 lkt1=-1.636594853e-07 wkt1=2.075371496e-08 pkt1=8.019445708e-14 kt2=-0.055045 at=3.067464233e+05 lat=-1.506450026e-1 ute=-1.385784630e-01 lute=1.721288918e-07 wute=2.098824955e-08 pute=-8.434453399e-14 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos lmin=1.5e-06 lmax=2e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.776540747e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=-2.549213958e-8 k1=0.64774 k2=-4.062982117e-02 wk2=-5.639589701e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.314351342e-09 wua=1.143930250e-16 ub=3.384790326e-18 wub=-1.259273157e-25 uc=2.287029360e-11 wuc=1.557672045e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.430616151e-03 wu0=3.611819316e-10 a0=2.344337631e+00 wa0=-3.209246786e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=6.288099588e-01 wags=-1.517505573e-7 b0=-3.213779458e-07 wb0=5.647731553e-14 b1=1.219520745e-07 wb1=3.906732134e-14 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-3.987916076e-01 wpclm=2.101588488e-7 pdiblc1=0.0 pdiblc2=5.861063403e-03 wpdiblc2=6.373713384e-10 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.807730911e-02 wdelta=-1.727429665e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.679973582e-01 wkt1=6.048039291e-8 kt2=-0.055045 at=232120.0 ute=-5.330936468e-02 wute=-2.079429080e-8 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos lmin=1e-06 lmax=1.5e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.809003889e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=4.930031285e-09 wvth0=-2.645654416e-09 pvth0=-3.469592893e-14 k1=0.64774 k2=-2.640731066e-02 lk2=-2.159908669e-08 wk2=1.054978798e-08 pk2=-2.458607936e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=3.563481218e+05 lvsat=-3.532211141e-01 wvsat=-8.373358456e-02 pvsat=1.271624269e-7 ua=-4.432672838e-09 lua=1.698344532e-15 wua=3.502116582e-16 pua=-3.581271464e-22 ub=5.077425525e-18 lub=-2.570528908e-24 wub=-6.194047604e-25 pub=7.494219887e-31 uc=-6.959988504e-11 luc=1.404302991e-16 wuc=4.253413536e-17 puc=-4.093901295e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=6.782934973e-04 lu0=1.142518560e-09 wu0=6.059998208e-11 pu0=4.564802806e-16 a0=4.265029687e+00 la0=-2.916868595e-06 wa0=-8.918103498e-07 pa0=8.669783791e-13 keta=-1.837780877e-02 lketa=8.804871275e-09 wketa=2.087257539e-09 pketa=-3.169824098e-15 a1=0.0 a2=0.46703705 ags=-8.394017210e-01 lags=2.229707009e-06 wags=4.170616793e-07 pags=-8.638295472e-13 b0=-1.845597958e-06 lb0=2.314764342e-12 wb0=7.638696298e-13 pb0=-1.074284875e-18 b1=-3.265632691e-07 lb1=6.811400691e-13 wb1=4.067744591e-15 pb1=5.315228222e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-3.987916076e-01 wpclm=2.101588488e-7 pdiblc1=0.0 pdiblc2=-4.316068790e-02 lpdiblc2=7.444712772e-08 wpdiblc2=1.165339136e-08 ppdiblc2=-1.672953388e-14 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.820286998e-02 ldelta=1.499586635e-08 wdelta=-3.690281126e-09 pdelta=2.980894185e-15 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.136865361e+00 lkt1=5.601832371e-07 wkt1=1.749616309e-07 pkt1=-1.738575045e-13 kt2=6.673269140e-03 lkt2=-9.372875802e-8 at=9.375863759e+05 lat=-1.071360039e+00 wat=-2.244009198e-01 pat=3.407875788e-7 ute=-1.725785291e-01 lute=1.811287128e-07 wute=4.189531444e-08 pute=-9.520388244e-14 ua1=3.961173043e-10 lua1=4.555550342e-16 wua1=1.199551055e-16 pua1=-1.821704207e-22 ub1=-4.331910094e-19 lub1=4.727740209e-25 wub1=1.246604198e-25 pub1=-1.893161698e-31 uc1=-9.137394491e-11 luc1=1.236381759e-16 wuc1=-6.162975822e-33 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos lmin=5e-07 lmax=1e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-1.383273890e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))' lvth0=-2.421681679e-07 wvth0=-1.280878447e-07 pvth0=9.308638543e-14 k1=0.64774 k2=4.671486150e-03 lk2=-5.325765846e-08 wk2=-4.157343061e-08 pk2=2.850949787e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.251798220e+05 lvsat=-1.177403696e-01 wvsat=-1.092638603e-02 pvsat=5.299701004e-8 ua=-2.744495711e-09 lua=-2.132553917e-17 wua=5.832544001e-17 pua=-6.079579086e-23 ub=2.147583121e-18 lub=4.139697062e-25 wub=1.689371852e-25 pub=-5.362647590e-32 uc=8.801917423e-11 luc=-2.012914367e-17 wuc=-4.587596908e-18 puc=7.061775235e-24 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.243084002e-04 lu0=1.604972749e-09 wu0=1.202097925e-09 pu0=-7.063123066e-16 a0=3.162376217e+00 la0=-1.793645124e-06 wa0=-8.243224845e-07 pa0=7.982315276e-13 keta=-9.734184308e-03 wketa=-1.024516416e-9 a1=0.0 a2=0.46703705 ags=1.232174113e+00 lags=1.194859274e-07 wags=-3.887201187e-07 pags=-4.301588976e-14 b0=1.641343734e-06 lb0=-1.237226247e-12 wb0=-7.479270759e-13 pb0=4.657143982e-19 b1=-5.977633844e-07 lb1=9.573994226e-13 wb1=5.032172473e-13 pb1=-4.553088544e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-7.494803984e-01 lpclm=3.572308902e-07 wpclm=3.819991618e-07 ppclm=-1.750459941e-13 pdiblc1=0.0 pdiblc2=-1.224731769e-01 lpdiblc2=1.552391912e-07 wpdiblc2=4.098440399e-08 ppdiblc2=-4.660771655e-14 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=8.955482801e-02 ldelta=-5.768716246e-08 wdelta=-3.009985496e-08 pdelta=2.988313861e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-4.634257031e-01 lkt1=-1.258194378e-07 wkt1=-3.895355686e-08 pkt1=4.404827111e-14 kt2=-0.085339 at=-2.611397998e+05 lat=1.497283734e-01 wat=1.874513112e-01 pat=-7.874775551e-8 ute=1.143924626e-01 lute=-1.111957227e-07 wute=-1.050540218e-07 pute=5.448679369e-14 ua1=8.848676004e-10 lua1=-4.231289869e-17 wua1=-7.923311778e-17 pua1=2.073365886e-23 ub1=8.392223872e-19 lub1=-8.233762476e-25 wub1=-3.632211689e-25 pub1=3.076668499e-31 uc1=3.0e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos lmin=3.5e-07 lmax=5e-07 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=-9.3275e-9 ll=0.0 lw=0.0 lwl=0.0 wint=2.9996e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.384395e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.384395e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.374095245e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-3.518222296e-08 wvth0=-4.691826920e-08 pvth0=5.098737924e-14 k1=0.64774 k2=-9.880974627e-02 lk2=4.134001423e-10 wk2=-7.209163233e-09 pk2=1.068629877e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-6.349913396e+05 lvsat=2.765262042e-01 wvsat=3.079660332e-01 pvsat=-1.123981376e-7 ua=-2.089620961e-09 lua=-3.609796024e-16 wua=-2.556599975e-16 pua=1.020543263e-22 ub=1.342280928e-18 lub=8.316437149e-25 wub=5.277782339e-25 pub=-2.397411800e-31 uc=8.329871954e-11 luc=-1.768085625e-17 wuc=4.642381736e-18 puc=2.274600662e-24 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.617178015e-03 lu0=-6.734110411e-10 wu0=-3.697947639e-10 pu0=1.089576960e-16 a0=-2.958862585e-01 wa0=7.147189353e-7 keta=-9.734184308e-03 wketa=-1.024516416e-9 a1=0.0 a2=0.46703705 ags=3.880677647e+00 lags=-1.254173673e-06 wags=-1.342202579e-06 pags=4.515125557e-13 b0=-2.572900751e-06 lb0=9.485127262e-13 wb0=5.186552042e-13 pb0=-1.912048343e-19 b1=4.315776363e-06 lb1=-1.591032535e-12 wb1=-1.295418087e-12 pb1=4.775623549e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.1819+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5373+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-6.071640265e-02 wpclm=4.449929380e-8 pdiblc1=0.0 pdiblc2=-9.474802234e-02 lpdiblc2=1.408594012e-07 wpdiblc2=-1.667449725e-09 ppdiblc2=-2.448611937e-14 pdiblcb=-0.025 drout=4.590528431e-01 wdrout=-1.180568585e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.262895256e-01 ldelta=-7.673979706e-08 wdelta=-4.803854818e-08 pdelta=3.918713155e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.742520936e-01 lkt1=8.725772376e-08 wkt1=1.589654272e-07 pkt1=-5.860339955e-14 kt2=-0.085339 at=6.923868878e+04 lat=-2.162408160e-02 wat=1.231653620e-01 pat=-4.540552651e-8 ute=1.761225950e-01 lute=-1.432123645e-7 ua1=1.000185802e-09 lua1=-1.021232603e-16 wua1=-1.357399589e-16 pua1=5.004121456e-23 ub1=-2.016054216e-18 lub1=6.575272393e-25 wub1=7.952024970e-25 pub1=-2.931553765e-31 uc1=3.0e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=-5.0625e-8 dwc=2.252e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.000816244375 mjs=0.3362 pbs=0.6587 cjsws=9.76976e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.5506845e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.ends sky130_fd_pr__pfet_01v8_lvt