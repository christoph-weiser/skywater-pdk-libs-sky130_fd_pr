* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8__toxe_mult=1.0
.param sky130_fd_pr__pfet_01v8__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8__overlap_mult=1.0
.param sky130_fd_pr__pfet_01v8__ajunction_mult=1.0
.param sky130_fd_pr__pfet_01v8__pjunction_mult=1.0
.param sky130_fd_pr__pfet_01v8__lint_diff=0.0
.param sky130_fd_pr__pfet_01v8__wint_diff=0.0
.param sky130_fd_pr__pfet_01v8__dlc_diff=0.0
.param sky130_fd_pr__pfet_01v8__dwc_diff=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_51=0.0
.include "sky130_fd_pr__pfet_01v8.pm3.spice"