* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_hvt__toxe_mult=0.948
.param sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_hvt__overlap_mult=0.91064
.param sky130_fd_pr__pfet_01v8_hvt__lint_diff=1.7325e-8
.param sky130_fd_pr__pfet_01v8_hvt__wint_diff=-3.2175e-8
.param sky130_fd_pr__pfet_01v8_hvt__dlc_diff=1.7325e-8
.param sky130_fd_pr__pfet_01v8_hvt__dwc_diff=-3.2175e-8
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=1.6702
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=-0.098011
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=0.00097522
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=6.9012e-20
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.00086508
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=-29674.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=-0.030352
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=1.8215e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=1.7209
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=-0.12703
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=-2.6856e-20
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=-0.0068783
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.00054806
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=-23641.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=-0.059296
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=1.9021e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=0.88917
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=-0.16742
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=0.22697
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=-0.05321
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=1.7862e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=-0.0030523
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0021726
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=0.02652
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=2.0425e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=-5.5786e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=0.56532
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=-0.11759
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=0.1273
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=-0.04025
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=5.1865e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=-0.0062951
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.0020197
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.036899
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=-6.1212e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=0.3705
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=-0.085417
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.18515
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=-0.063572
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=4.5105e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=-0.0087946
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.0016238
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=0.029425
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=3.4914e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=0.58901
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=-0.052472
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=0.051784
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=-0.063375
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=4.024e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=-0.010302
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.0021038
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=0.025149
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=4.112e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=2.3478
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=-0.15288
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=-1.3862e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=-0.013041
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0015364
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=-27670.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=-0.053351
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=0.0010756
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=3.3792e-19
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=-15990.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=-0.059438
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=1.0152e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=1.0669
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=-0.11315
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=0.013182
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=0.0065099
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=0.0021339
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=3.4578e-19
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=-29944.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=0.037342
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=4.1649e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=1.2977
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=-0.045339
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=-0.073336
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=-0.012277
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0045307
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=4.1908e-20
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=-10537.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.045267
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=7.7724e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=1.4783
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=7.2706e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=-0.071099
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=-0.0037068
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=0.00973
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=0.2504
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.0023319
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.020152
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=-0.010112
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=-1.437e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=-1.3981e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=9.452e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=-0.10271
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=0.025822
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=-0.010134
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=-0.17771
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.0035013
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=0.013621
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=-0.011751
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=-0.010705
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=-1.7178e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=1.079e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=-0.067375
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=0.067597
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=-0.042239
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=0.27193
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.0041731
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=-0.017373
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=0.27144
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=0.0048327
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=0.00227
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=-0.00843
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=-3.3818e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=1.4661e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=-0.066337
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=0.037844
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=-0.021169
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=-24444.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=1.2545
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.00041791
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=-0.049892
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=-0.0042041
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=9.4745e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=4.124e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=-0.12375
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=-6505.6
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=0.66146
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.00089379
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=-0.071254
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=-8.1586e-5
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=1.6305e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=1.0152e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=-0.093754
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=-28762.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=0.70713
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.0012256
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=-0.001682
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0028259
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=1.3012e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=2.539e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=-0.04469
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=0.52823
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=0.0026198
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=13859.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.016554
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=-0.006883
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=1.1056e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=5.0826e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=-0.073286
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=-0.008952
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=0.011728
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=0.28249
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0023179
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=0.016121
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=-0.011899
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=-1.6357e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=7.6564e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=-0.06502
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=-0.077046
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.038942
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=-0.039498
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=0.12738
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0031187
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=0.0029058
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=-0.0081995
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=-2.5441e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=1.0061e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=-0.066055
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.016281
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=-0.015815
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=0.26745
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.0046376
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=0.0014783
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=-0.0077373
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=-3.3629e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=1.4023e-18
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=1.3543e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=-0.04378
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=-0.038207
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=-0.044188
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=0.36554
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=0.0039903
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.01708
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=-0.0066951
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=-4.1477e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=1.324e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=-4.5976e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=-0.084594
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=-26795.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=1.0827
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=0.00042769
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=-0.071575
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=0.00045233
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=0.0076182
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=1.5074e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=7.5942e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=-0.048212
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=-20619.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=0.71624
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.00066193
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=-0.050276
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=0.31532
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.00084832
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=-0.0077162
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=0.001811
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=-2.852e-13
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=3.5019e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=-0.050657
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=-11016.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=-2879.9
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=0.28888
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=0.00033371
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.028527
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=-0.0086212
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=-1.3033e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=1.7081e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=-0.056202
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=0.11511
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0033142
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=0.0065868
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=-0.0096254
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=-2.915e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=1.086e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=-0.066547
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.017504
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=-0.021718
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=-0.025453
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.004512
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=0.0029878
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=-0.010442
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=-3.7793e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=1.4138e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=-0.058137
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.045741
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=-0.048361
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=0.36762
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0049774
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.017746
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=-0.0066393
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=-4.132e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=1.5608e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=-0.045427
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=-0.0082778
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=0.0056012
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=-0.00067009
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=0.0017417
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=0.97578
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0092277
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.008761
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=-0.011014
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=-5.3257e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=1.8573e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=-0.034623
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=-0.088188
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=-18897.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=1.1748
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.00083903
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=-0.073728
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=-0.019298
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=2.86e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=-1.7396e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=-0.086699
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=-4248.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=0.42507
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=0.00024638
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=-0.085301
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=0.0015551
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=-1.6895e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=1.885e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=2.5238e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=-0.06692
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=-11755.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=0.35759
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.00068645
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=-0.0035656
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=8.2421e-5
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=2.8428e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=1.9174e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=1.8e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=-0.047344
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=-32711.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=0.97073
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0021523
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=0.013441
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=-0.0091659
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=-0.011769
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=-1.0721e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=1.3365e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=-0.12761
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=7.2095e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=5.0779e-8
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=1.0947
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0050028
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=0.046227
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=0.49911
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.003451
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=-0.0087503
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=-0.017093
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=-1.9758e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=9.821e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=-0.094876
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=-1.0283e-7
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=2.3178e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=0.69604
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=0.0062132
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=0.013867
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=-0.018297
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=6.1158e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=1.2575e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=-0.099857
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=5.6678e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=1.5052e-8
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=-1.0273e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=0.74962
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0031442
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=0.033856
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=-0.012048
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=1.0374e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=4.574e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=-0.076379
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=9.5235e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=1.91e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=-2.6206e-7
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=0.5372
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.0060424
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=0.0034632
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=-0.016469
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=7.736e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=3.488e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=-0.087212
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=2.2787
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.0025449
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=-50000.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.040102
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=-0.0018016
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=5.933e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=2.2929e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=-0.19968
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=-45149.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=1.9521
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=0.0021813
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.00501
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=-0.0085993
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=5.5697e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=6.3421e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=-0.19674
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=-0.093014
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=-38889.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=1.6445
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.0057123
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.091479
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=-0.023719
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=4.3063e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=8.5174e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=-0.08843
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=1.0665e-7
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=9.4459e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=1.3174
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0047
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=0.034666
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=-0.014806
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=7.2762e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=-4.3961e-20
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=2.8498e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=-0.061848
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=1.1443e-7
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=-1.6295e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=0.73413
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.003296
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=0.041686
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=-0.0061916
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=2.8632e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=-4.6452e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=5.5996e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=-0.069356
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=9.4887e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=2.3137e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=0.4916
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0024626
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=0.03279
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=-0.0078584
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=-0.0088326
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=-1.474e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=5.7719e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=-0.067651
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=7.7369e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=7.0231e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=0.3621
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=0.0019517
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.026283
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=2.0889
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.0012322
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=-0.039462
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=-0.016442
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=2.1814e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=1.5922e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=-0.13831
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=-40582.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=-50000.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=3.6882
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.015631
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.074708
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=-0.0080946
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=2.0e-9
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=1.1367e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=-0.075714
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=-24472.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=2.5262
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=0.0012175
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=-0.023234
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=-0.007354
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=2.5998e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=1.7343e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=-0.19561
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=-30755.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=1.8113
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.001795
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=-0.012419
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=-0.0068842
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=5.2165e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=-1.2533e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=-0.15886
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=-29893.59829279
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.00124944
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=1.72013046
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=-0.04127798
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.0010617
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=3.46701e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=1.396e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=-0.103349
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=-14190.02188706
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=3.06099e-5
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.96707997
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=-0.07541995
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.00703588
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=5.6917e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=-2.9419e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=-0.082426
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=-0.072042
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=-7.6647e-8
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=-26609.98832683
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=0.0003282
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=1.21669943
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=-0.05314867
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.012422
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=6.42999e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=1.03621e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=-0.09478604
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=-16214.19463122
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=-0.00051934
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=1.11233043
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=-0.071217
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.00941368
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=-1.5565e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=2.02164e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=-2.0137e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=-0.109857
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=-24608.56214497
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=0.00160218
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=0.39679982
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=-0.06057999
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=0.00330583
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=5.29585e-10
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=1.77615e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=-1.065e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=-0.036074
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=-39429.59956441
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=0.00036125
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=0.53532009
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=-0.0623438
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.01331141
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=-0.0066348
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=-30180.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=-0.001025
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.08346
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=-0.00056441
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=0.0086191
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=0.0054426
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=-37723.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=-30636.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=-0.00052667
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=-0.00043348
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=0.0051619
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=-27201.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.00143932
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=0.0013145
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=1.243108
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=-0.044733
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=-0.005647
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=4.11678e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=-6.27298e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=-0.00026826
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=-0.00136297
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=-0.10590279
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=4.2886e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=-7.09239e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=-7.29796e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=-25393.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=0.0012886
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.00148104
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=0.90432662
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=-0.05008
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=-0.0047585
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=4.5847e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=-1.17829e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=-0.00027604
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=-0.10757491
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=-0.00140248
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=4.41291e-12
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=3.018e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=-4.9911e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=-23783.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.00101288
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=0.0013326
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=0.66438835
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=-0.052569
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=-0.0044981
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=4.91938e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=-1.57174e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=-0.00018878
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=-0.10868729
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=-0.00095916
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=1.34608e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=-2.22611e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=-21900.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.00045176
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=0.0013726
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=0.49989482
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=-0.054622
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=-0.0029267
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=5.1504e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=-1.84303e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=-8.42008e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=-0.10941523
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=-0.0004278
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=-0.0004278
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=-0.10941523
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=1.34608e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=-2.22613e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=-23535.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.00045176
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=0.0015171
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=0.49989469
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=-0.034774
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=-0.013873
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=5.1504e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=-1.84303e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=-8.42007e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=-0.0001157
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=-434810.89830208
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=-0.00046359
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.00047433
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=-0.0245589
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=1.562e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=3.46622e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=-19223.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=0.0022188
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=0.81033175
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=0.019208
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=0.0049685
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=2.61701e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=3.89042e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=-15187.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=-0.00058999
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.046929
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=-0.0016053
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=4.61965e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=-1.56897e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.00031999
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=-0.10432908
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=-4.53896e-13
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=1.91787e-6
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=-18965.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=2.59995e-5
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=0.0012435
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=0.51671158
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=-0.056768
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=-0.0024326
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=-0.0012624
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=2.20238e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=1.67256e-21
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=7.9727e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.00057533
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=-0.08465745
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=-8.16075e-13
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=3.44709e-6
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=-17711.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=4.67463e-5
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=0.00053342
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=0.94327401
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=-0.047237
.include "sky130_fd_pr__pfet_01v8_hvt__fs.pm3.spice"