* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.model sky130_fd_pr__diode_pw2nd_11v0__no_rs d level=3.0 tlevc=1.0 area=1.0e+12 cj='0.0008512*1e-12*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult' mj=0.295 pb=0.72468 cjsw='8.5204e-011*1e-6*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult' mjsw=0.037586 php=0.29067 cta=0.00067434 ctp=0.0002493 tpb=0.001344 tphp=0.00099005 js=3.75e-016 jsw=5.84e-017 n=1.0773 rs=0 ik='1.3e-009/1e-12' ikr='0/1e-12' vb=12.636 ibv=0.00106 trs=0 eg=0.92 xti=0.76 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0