* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_b__toxe_mult=1.0365
.param sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult=1.2
.param sky130_fd_pr__rf_nfet_01v8_b__overlap_mult=0.98
.param sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult=1.1505
.param sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult=1.1793
.param sky130_fd_pr__rf_nfet_01v8_b__lint_diff=-1.21275e-8
.param sky130_fd_pr__rf_nfet_01v8_b__wint_diff=2.252e-8
.param sky130_fd_pr__rf_nfet_01v8_b__rshg_diff=7.0
.param sky130_fd_pr__rf_nfet_01v8_b__dlc_diff=-11.107e-9
.param sky130_fd_pr__rf_nfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_b__xgw_diff=4.504e-8
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_0=0.016061
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_0=7256.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_0=0.0079631
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_0=-0.0019138
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_1=0.020817
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_1=9830.4
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_1=0.014994
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_1=-0.002237
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_2=0.0086842
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_2=19450.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_2=0.032627
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_2=-0.0030221
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_3=0.025003
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_3=1653.2
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_3=0.0026575
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_3=-0.0083307
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_4=0.00020419
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_4=12334.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_4=0.015143
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_4=-0.0053582
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_5=0.0016884
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_5=11246.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_5=0.034079
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_5=-0.0028787
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_6=-0.006203
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_6=0.0065467
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_6=-4610.9
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_6=0.001022
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_7=0.013198
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_7=-0.0055047
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_7=-0.0028156
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_7=9383.7
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_8=0.031946
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_8=-0.0050561
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_8=-0.0043506
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_8=12165.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_0=0.0068964
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_0=-0.0035814
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_0=0.040659
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_0=-2843.6
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_1=0.019365
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_1=-0.0039029
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_1=0.0080414
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_1=11376.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_2=0.035011
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_2=-0.0035828
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_2=0.0072093
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_2=24875.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_3=526.28
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_3=0.0028165
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_3=-0.0086312
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_3=0.018526
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_4=14947.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_4=0.017688
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_4=-0.008178
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_4=-0.0046622
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_5=40210.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_5=0.035635
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_5=-0.0070625
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_5=-0.0049699
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_6=-4885.3
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_6=0.0013795
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_6=-0.0060867
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_6=0.0069395
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_7=-0.0068351
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_7=3065.3
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_7=0.016371
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_7=-0.012469
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_8=-0.0078852
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_8=-0.0064297
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_8=34241.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_8=0.033541
.include "sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"