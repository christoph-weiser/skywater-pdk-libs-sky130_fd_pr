* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.include "../../models/parasitics/sky130_fd_pr__model__parasitic__diode_pw2dn__extended_drain.model.spice"
.include "../diode_pw2nd_05v5/sky130_fd_pr__diode_pw2nd_05v5__extended_drain.model.spice"
.subckt sky130_fd_pr__nfet_20v0 d g s b w=60u l=2u m=1 t=30 ad=0 as=0 pd=0 ps=0 nrd=2 nrs=2 mf=1 sa=0 sb=0
.param rdrift_tnom=1.934600e+004
.param vgdep_tnom=6.000000e-002
.param vth_tnom=7.000000e-001
.param vbdep_tnom=-1.224000
.param vth2=+1.048000e-001
.param hvvsat_tnom=3.893600
.param avsat_tnom=9.407600e-001
.param deltaw=9.000000e-001
.param hvnel_n20vhv1=2.95
.param hvvbdep=-2.490600e-002
.param sky130_fd_pr__nfet_20v0__vgdep_mult=1
.param n20vhv1res_vth0_diff=0.0
.param sky130_fd_pr__nfet_20v0__vbdep_mult=1
.param sky130_fd_pr__nfet_20v0__avsat_mult=1
.param sky130_fd_pr__nfet_20v0__pgatejunction_mult=4.6689e-1
.param sky130_fd_pr__nfet_20v0__mjswgatejunction_mult=1.0
.param sky130_fd_pr__nfet_20v0__pbswgatejunction_mult=1.0
.param w_n20vhv1=29.41
.param nrd_n20vhv1=2.0
.param nrs_n20vhv1=2.0
.param ad_n20vhv1='294.5*0.5'
.param as_n20vhv1=8.7
.param pd_n20vhv1='91.5*0.5'
.param ps_n20vhv1=60.58
.param delvto_n20vhv1=0.0
.param tc1_rdrift=0.00671814786081909
.param tc1_vgdep=0.00067352380952381
.param tc1_vth=0.00573669467787115
.param tc1_vbdep=-0.000337318979879533
.param tc1_hvvsat=0.0070429485950945
.param tc1_avsat=0.00120508503584265
.param tc2_rdrift=1.77312980397369e-05
.param tc2_vgdep=7.92380952380953e-06
.param tc2_vth=-0.000036750700280112
.param tc2_vbdep=-1.67576573112905e-05
.param tc2_hvvsat=-6.16729946550226e-06
.param tc2_avsat=-1.16883863966948e-05
.param rdrift='rdrift_tnom*((w_n20vhv1-deltaw)/w_n20vhv1)*(1+tc1_rdrift*(temper-30)+tc2_rdrift*(temper-30)*(temper-30))*sky130_fd_pr__nfet_20v0__rdrift_mult'
.param vgdep='vgdep_tnom*(1+tc1_vgdep*(temper-30)+tc2_vgdep*(temper-30)*(temper-30))*sky130_fd_pr__nfet_20v0__vgdep_mult'
.param vth='vth_tnom*(1+tc1_vth*(temper-30)+tc2_vth*(temper-30)*(temper-30))+n20vhv1res_vth0_diff'
.param vbdep='vbdep_tnom*(1+tc1_vbdep*(temper-30)+tc2_vbdep*(temper-30)*(temper-30))*sky130_fd_pr__nfet_20v0__vbdep_mult'
.param hvvsat='hvvsat_tnom*(1+tc1_hvvsat*(temper-30)+tc2_hvvsat*(temper-30)*(temper-30))*sky130_fd_pr__nfet_20v0__hvvsat_mult'
.param avsat='avsat_tnom*(1+tc1_avsat*(temper-30)+tc2_avsat*(temper-30)*(temper-30))*sky130_fd_pr__nfet_20v0__avsat_mult'
m1 d1 g s b sky130_fd_pr__nfet_20v0__base w=w_n20vhv1 l=hvnel_n20vhv1 ad=0 as=0 pd=0 ps=0 nrd=nrd_n20vhv1 nrs=nrs_n20vhv1 delvto=delvto_n20vhv1 m=m
rldd d d1 r='abs((1/w_n20vhv1)*(rdrift/(1+vgdep*(v(g,s)-vth-vbdep*v(b,s))))*(1+pwr((abs(v(d,s)+vth2-min(v(d1,s),60))/(hvvsat*(1+hvvbdep*v(b,s)))),avsat)))' tc1=0 tc2=0 m='m'
dndrain1 b d sky130_fd_pr__model__parasitic__diode_ps2dn__extended_drain area='0.5*ad_n20vhv1' pj='0.5*pd_n20vhv1' m=m
dndrain2 b d1 sky130_fd_pr__model__parasitic__diode_ps2dn__extended_drain area='0.5*ad_n20vhv1' pj='0.5*pd_n20vhv1' m=m
dnsrc b s sky130_fd_pr__diode_pw2nd_05v5__extended_drain area='as_n20vhv1' pj='ps_n20vhv1-w_n20vhv1' m=m
.model sky130_fd_pr__nfet_20v0__base.0 nmos lmin=4.95e-07 lmax=3.05e-06 wmin=1.9995e-05 wmax=6.0005e-5 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.6507e-08+sky130_fd_pr__nfet_20v0__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.1346e-08+sky130_fd_pr__nfet_20v0__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.1292e-9 dwb=-1.6944e-9 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__nfet_20v0__toxe_mult' dtox=0.0 ndep=1.7e+17 nsd=1.0e+20 rshg=0.1 rsh='1.0*sky130_fd_pr__nfet_20v0__rshn_mult' vth0='0.80788+sky130_fd_pr__nfet_20v0__vth0_diff' k1=0.88325 k2='-0.022723+sky130_fd_pr__nfet_20v0__k2_diff' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.19251 dvt0w=0.16 dvt1w=6909100.0 dvt2w=-0.036016 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.1160e+5 ua=-1.321700e-10 ub=9.6801e-19 uc=1.0857e-10 rdsw=724.62 prwb=0.05626 prwg=0.048 wr=1.0 u0=0.17559 a0=2.1951 keta=-0.01066 a1=0.0 a2=0.65972622 ags=0.18589 b0=3.2933e-8 b1=0.0 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff=-0.20613 nfactor=0.2786 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.056336 etab=-0.01932 dsub=0.504 voffl=-4.2579486e-7 minv=0.0 pclm=1.2848 pdiblc1=0.21098 pdiblc2=0.0002 pdiblcb=-0.26831 drout=0.36075 pscbe1=2.2576e+9 pscbe2=1.68e-6 pvag=1.99 delta=0.0246 alpha0=9.8435e-9 alpha1=0.0 beta0=36.96 fprout=10.125 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-16 bgidl=1058000000.0 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1=-0.35073 kt2=-0.019151 at=49600.0 ute=-1.2986 ua1=3.0044e-9 ub1=-3.4025e-18 uc1=-5.9821e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1000000e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.0773 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.636 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.00099005 tpbswg=0.0 tcj=0.00067434 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.90e-010*sky130_fd_pr__nfet_20v0__overlap_mult' cgso='2.90e-010*sky130_fd_pr__nfet_20v0__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-011*sky130_fd_pr__nfet_20v0__overlap_mult' cgdl='5e-011*sky130_fd_pr__nfet_20v0__overlap_mult' cf=0.0 clc=1.0e-7 cle=0.6 dlc='7.20e-07+sky130_fd_pr__nfet_20v0__dlc_diff' dwc='0.0+sky130_fd_pr__nfet_20v0__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=4.0 voffcv=-0.4104 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0008512*sky130_fd_pr__nfet_20v0__ajunction_mult' mjs=0.295 pbs=0.72468 cjsws='8.5204e-011*sky130_fd_pr__nfet_20v0__pjunction_mult' mjsws=0.037586 pbsws=0.29067 cjswgs='5.4e-011*sky130_fd_pr__nfet_20v0__pgatejunction_mult*sky130_fd_pr__nfet_20v0__pjunction_mult' mjswgs='0.78692*sky130_fd_pr__nfet_20v0__mjswgatejunction_mult' pbswgs='0.54958*sky130_fd_pr__nfet_20v0__pbswgatejunction_mult' saref=1.81e-6 sbref=1.81e-6 wlod=0.0 kvth0=1.1e-8 lkvth0=0.0 wkvth0=6.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-4.5e-8 lku0=0.0 wku0=2.0e-7 pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.3 steta0=0.0 tku0=0.0
.ends sky130_fd_pr__nfet_20v0