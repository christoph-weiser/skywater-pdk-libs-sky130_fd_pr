* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre=0.0
.subckt sky130_fd_pr__nfet_01v8 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__nfet_01v8__model.0 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.540388+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.031308211 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.2609486+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.68119 eta0=0.08 etab=-0.07 u0=0.0325965 ua=-7.5800507e-10 ub=1.7355048e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.278231 ags=0.455362 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.00096922 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.1 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.540388+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.031308211 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.2609486+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.68119 eta0=0.08 etab=-0.07 u0=0.0325965 ua=-7.5800507e-10 ub=1.7355048e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.278231 ags=0.455362 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.00096922 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.2 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.410417073e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-5.191407026e-09 wvth0=-6.538421294e-08 pvth0=5.192478117e-13 k1=5.415461066e-01 lk1=-5.403836471e-09 wk1=-6.805969803e-08 pk1=5.404951391e-13 k2=-3.188143178e-02 lk2=4.552224783e-09 wk2=5.733390449e-08 pk2=-4.553163998e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.611814635e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.849282207e-09 wvoff=2.329115422e-08 pvoff=-1.849663751e-13 nfactor=2.681509861e+00 lnfactor=-2.540174125e-09 wnfactor=-3.199273050e-08 pnfactor=2.540698214e-13 eta0=0.08 etab=-0.07 u0=3.259529717e-02 lu0=9.552236187e-12 wu0=1.203075470e-10 pu0=-9.554207004e-16 ua=-7.576149024e-10 lua=-3.098510305e-18 wua=-3.902480707e-17 pua=3.099149590e-22 ub=1.736245703e-18 lub=-5.883870307e-27 wub=-7.410558008e-26 pub=5.885084267e-31 uc=4.876986983e-11 luc=3.749415156e-18 wuc=4.722275825e-17 puc=-3.750188736e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.270180686e+00 la0=6.393145682e-08 wa0=8.051975054e-07 pa0=-6.394464716e-12 ags=4.563758116e-01 lags=-8.051170500e-09 wags=-1.014020754e-07 pags=8.052831618e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=1.950584888e-24 lb1=1.244887590e-30 wb1=1.567898546e-29 pb1=-1.245144435e-34 keta=-8.287828103e-03 lketa=-4.024521921e-09 wketa=-5.068764537e-08 pketa=4.025352261e-13 dwg=0.0 dwb=0.0 pclm=6.802472480e-02 lpclm=-3.312292541e-07 wpclm=-4.171733015e-06 ppclm=3.312975933e-11 pdiblc1=0.39 pdiblc2=3.074732737e-03 lpdiblc2=-1.011774984e-11 wpdiblc2=-1.274300217e-10 ppdiblc2=1.011983733e-15 pdiblcb=-0.025 drout=0.56 pscbe1=7.580457839e+08 lpscbe1=-2.677570371e+01 wpscbe1=-3.372319497e+02 ppscbe1=2.678122808e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.131869552e-01 lkt1=1.246457536e-09 wkt1=1.569875846e-08 pkt1=-1.246714705e-13 kt2=-4.539675534e-02 lkt2=6.624655971e-10 wkt2=8.343555311e-09 pkt2=-6.626022770e-14 at=140000.0 ute=-1.816360577e+00 lute=2.351137911e-08 wute=2.961187614e-07 pute=-2.351622998e-12 ua1=3.613688642e-10 lua1=1.163517897e-16 wua1=1.465415860e-15 pua1=-1.163757954e-20 ub1=-6.204394793e-19 lub1=-1.523218368e-25 wub1=-1.918447805e-24 pub1=1.523532638e-29 uc1=1.691037604e-11 luc1=-8.582070437e-18 wuc1=-1.080886007e-16 puc1=8.583841090e-22 kt1l=0.0 prt=0.0 tvoff=9.565096041e-04 ltvoff=1.009394309e-10 wtvoff=1.271301828e-09 ptvoff=-1.009602567e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.3 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.312943148e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.322780398e-08 wvth0=5.629118589e-08 pvth0=3.966593064e-14 k1=5.306153844e-01 lk1=3.767945204e-08 wk1=1.370579661e-07 pk1=-2.679732626e-13 k2=-2.280303039e-02 lk2=-3.123016719e-08 wk2=-1.024852280e-07 pk2=1.746084733e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.380153891e-01 ldsub=8.665203596e-08 wdsub=2.198914673e-06 pdsub=-8.666991401e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.574732096e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.276674851e-08 wvoff=-4.366083040e-08 pvoff=7.892393489e-14 nfactor=2.685068065e+00 lnfactor=-1.656478334e-08 wnfactor=-8.053921037e-07 pnfactor=3.302412623e-12 eta0=7.417407812e-02 leta0=2.296278953e-08 weta0=5.827123885e-07 peta0=-2.296752721e-12 etab=-6.490694912e-02 letab=-2.007418872e-08 wetab=-5.094101673e-07 petab=2.007833043e-12 u0=3.248454674e-02 lu0=4.460735132e-10 wu0=1.276765103e-08 pu0=-5.080474799e-14 ua=-7.764702823e-10 lua=7.121970541e-17 wua=1.337627886e-15 pua=-5.116142358e-21 ub=1.732606123e-18 lub=8.461481542e-27 wub=-6.771514625e-25 pub=2.965405330e-30 uc=5.865001446e-11 luc=-3.519303660e-17 wuc=-3.247378503e-16 puc=1.091058657e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.394640551e+00 la0=-4.266253605e-07 wa0=-1.135517398e-06 pa0=1.254835905e-12 ags=4.565489758e-01 lags=-8.733694935e-09 wags=-1.442020674e-06 pags=6.089312598e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=4.466545308e-24 lb1=-8.671735184e-30 wb1=-3.135797092e-29 pb1=6.088106153e-35 keta=-1.628561723e-02 lketa=2.749865195e-08 wketa=8.778174682e-08 pketa=-1.432399447e-13 dwg=0.0 dwb=0.0 pclm=-6.034433030e-01 lpclm=2.315352577e-06 wpclm=8.547745203e-06 ppclm=-1.700388599e-11 pdiblc1=0.39 pdiblc2=3.180469299e-03 lpdiblc2=-4.268769279e-10 wpdiblc2=-1.236623145e-08 ppdiblc2=4.925104822e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.039311704e+08 lpscbe1=1.865162878e+02 wpscbe1=6.744638995e+02 ppscbe1=-1.309462218e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.113156351e-01 lkt1=-6.129324575e-09 wkt1=3.339716880e-08 pkt1=-1.944295071e-13 kt2=-4.405890304e-02 lkt2=-4.610660505e-09 wkt2=-1.658575532e-08 pkt2=3.199830113e-14 at=1.381635522e+05 lat=7.238333404e-03 wat=1.836826724e-01 pat=-7.239826817e-7 ute=-1.758708369e+00 lute=-2.037239891e-07 wute=-1.605937187e-06 pute=5.145303895e-12 ua1=6.189646349e-10 lua1=-8.989583341e-16 wua1=-5.175777008e-15 pua1=1.453858917e-20 ub1=-9.417373089e-19 lub1=1.114069061e-24 wub1=5.182191606e-24 pub1=-1.275174445e-29 uc1=1.117151042e-14 luc1=5.802590764e-17 wuc1=1.716226603e-16 puc1=-2.440939101e-22 kt1l=0.0 prt=0.0 tvoff=1.141105832e-03 ltvoff=-6.266440175e-10 wtvoff=-6.016216739e-10 ptvoff=-2.713923907e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.4 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.494174425e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.957994842e-09 wvth0=-2.414923493e-08 pvth0=1.958398815e-13 k1=5.524216916e-01 lk1=-4.657188206e-09 wk1=-2.408938554e-07 pk1=4.658149077e-13 k2=-3.958824177e-02 lk2=1.358085705e-09 wk2=5.741552014e-08 pk2=-1.358365905e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.826472000e-01 wdsub=-2.265187257e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.646821291e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.229267677e-09 wvoff=6.031935016e-08 pvoff=-1.229521299e-13 nfactor=2.678822107e+00 lnfactor=-4.438343342e-09 wnfactor=6.669268918e-07 pnfactor=4.439259061e-13 eta0=8.614587586e-02 leta0=-2.802881704e-10 weta0=-6.147143873e-07 peta0=2.803459994e-14 etab=-7.523317378e-02 letab=-2.596811357e-11 wetab=5.234253492e-07 petab=2.597347131e-15 u0=3.237751711e-02 lu0=6.538700426e-10 wu0=2.028547342e-08 pu0=-6.540049491e-14 ua=-7.764744977e-10 lua=7.122788960e-17 wua=2.371947050e-15 pua=-7.124258534e-21 ub=1.767483152e-18 lub=-5.925178081e-26 wub=-2.202269457e-24 pub=5.926400564e-30 uc=3.956786110e-11 luc=1.854697008e-18 wuc=3.327825359e-16 puc=-1.855079669e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.144279014e+04 lvsat=-2.801156853e-03 wvsat=-1.443087814e-01 pvsat=2.801734788e-7 a0=1.168136717e+00 la0=1.312866340e-08 wa0=1.871669356e-07 pa0=-1.313137211e-12 ags=4.711814167e-01 lags=-3.714237396e-08 wags=-2.190868585e-07 pags=3.715003717e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.737729786e-03 lketa=8.961562150e-09 wketa=4.756811009e-07 pketa=-8.963411100e-13 dwg=0.0 dwb=0.0 pclm=5.772212616e-01 lpclm=2.310885410e-08 wpclm=9.800760065e-07 ppclm=-2.311362192e-12 pdiblc1=4.125418191e-01 lpdiblc1=-4.376462613e-08 wpdiblc1=-2.254646989e-06 ppdiblc1=4.377365565e-12 pdiblc2=2.903662834e-03 lpdiblc2=1.105389482e-10 wpdiblc2=1.869617316e-08 ppdiblc2=-1.105617546e-14 pdiblcb=-2.323678196e-02 lpdiblcb=-3.423263134e-09 wpdiblcb=-1.763581824e-07 ppdiblcb=3.423969421e-13 drout=5.386779783e-01 ldrout=4.139640670e-08 wdrout=2.132642090e-06 pdrout=-4.140494760e-12 pscbe1=7.616967335e+08 lpscbe1=7.436525565e+01 wpscbe1=3.831116922e+03 ppscbe1=-7.438059869e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.155015891e-07 lalpha0=-3.601487383e-13 walpha0=-1.855398618e-11 palpha0=3.602230442e-17 alpha1=8.524164958e-01 lalpha1=-4.691592759e-09 walpha1=-2.416994369e-07 palpha1=4.692560729e-13 beta0=1.405701548e+01 lbeta0=-3.825027979e-07 wbeta0=-1.970561291e-05 pbeta0=3.825817159e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.108273075e-01 lkt1=-7.077405665e-09 wkt1=-4.313582271e-07 pkt1=7.078865876e-13 kt2=-4.500785316e-02 lkt2=-2.768287140e-09 wkt2=-1.427198239e-07 pkt2=2.768858293e-13 at=1.382262563e+05 lat=7.116594264e-03 wat=1.774109683e-01 pat=-7.118062559e-7 ute=-1.804785838e+00 lute=-1.142652292e-07 wute=-4.842415092e-06 pute=1.142888044e-11 ua1=2.781043722e-10 lua1=-2.371829062e-16 wua1=-9.906480707e-15 pua1=2.372318418e-20 ub1=-4.320543041e-19 lub1=1.245266422e-25 wub1=5.029467871e-24 pub1=-1.245523345e-29 uc1=3.127958242e-11 luc1=-2.681274377e-18 wuc1=-9.223536801e-17 puc1=2.681827578e-22 kt1l=0.0 prt=0.0 tvoff=8.330500355e-04 ltvoff=-2.855800110e-11 wtvoff=-3.470719482e-09 ptvoff=2.856389319e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.5 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.381666099e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.634506540e-09 wvth0=2.037931952e-07 pvth0=-1.876472530e-14 k1=5.410715732e-01 lk1=6.028789400e-09 wk1=9.056609530e-07 pk1=-6.136503927e-13 k2=-3.396882486e-02 lk2=-3.932516640e-09 wk2=-3.578547329e-07 pk2=2.551345389e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.765676518e-01 ldsub=-2.767219905e-07 wdsub=-5.168671357e-06 pdsub=2.733589631e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.636399368e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.480582220e-10 wvoff=-8.720622728e-09 pvoff=-5.795196202e-14 nfactor=2.556416381e+00 lnfactor=1.108049336e-07 wnfactor=2.434933257e-06 pnfactor=-1.220627335e-12 eta0=1.938363928e-01 leta0=-1.016694022e-07 weta0=-4.364912258e-06 peta0=3.558793393e-12 etab=-1.412592556e-01 letab=6.213666359e-08 wetab=9.895353030e-07 petab=-4.362386488e-13 u0=3.454453944e-02 lu0=-1.386351145e-09 wu0=-3.972544891e-08 pu0=-8.901051683e-15 ua=-5.483446588e-10 lua=-1.435531599e-16 wua=-5.269140955e-15 pua=6.971884766e-23 ub=1.596618779e-18 lub=1.016146341e-25 wub=4.942935509e-24 pub=-8.007098789e-31 uc=1.315963194e-11 luc=2.671767505e-17 wuc=1.993682048e-16 puc=-5.990024203e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.905634652e+04 lvsat=-5.543536001e-04 wvsat=9.438481717e-02 pvsat=5.544679744e-8 a0=1.276262256e+00 la0=-8.867001772e-08 wa0=-4.905838533e-06 pa0=3.481856136e-12 ags=2.377884906e-01 lags=1.825937985e-07 wags=3.306599856e-06 pags=3.956190354e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.567290278e-03 lketa=-7.404699696e-10 wketa=-7.188215256e-07 pketa=2.282663898e-13 dwg=0.0 dwb=0.0 pclm=6.378922917e-01 lpclm=-3.401207138e-08 wpclm=-2.626928087e-06 ppclm=1.084581664e-12 pdiblc1=3.855766103e-01 lpdiblc1=-1.837725957e-08 wpdiblc1=4.424302360e-07 ppdiblc1=1.838105116e-12 pdiblc2=1.346831978e-03 lpdiblc2=1.576273404e-09 wpdiblc2=2.234040849e-08 ppdiblc2=-1.448717200e-14 pdiblcb=-2.852643607e-02 lpdiblcb=1.556872156e-09 wpdiblcb=3.527163648e-07 ppdiblcb=-1.557193370e-13 drout=5.985615139e-01 ldrout=-1.498310375e-08 wdrout=-3.856946992e-06 pdrout=1.498619506e-12 pscbe1=8.606637269e+08 lpscbe1=-1.881078310e+01 wpscbe1=-6.067624304e+03 ppscbe1=1.881466414e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.693400696e-08 lalpha0=-2.108595796e-13 walpha0=-2.693956398e-12 palpha0=2.109030842e-17 alpha1=8.451670084e-01 lalpha1=2.133698127e-09 walpha1=4.833988737e-07 palpha1=-2.134138352e-13 beta0=1.379525039e+01 lbeta0=-1.360546335e-07 wbeta0=6.476296493e-06 pbeta0=1.360827043e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.102204899e-01 lkt1=-7.648715918e-09 wkt1=2.886557859e-07 pkt1=3.000347447e-14 kt2=-4.858103395e-02 lkt2=5.958125495e-10 wkt2=2.158932027e-07 pkt2=-6.074331455e-14 at=1.689204043e+05 lat=-2.178151638e-02 wat=-6.794527531e-01 pat=9.491894162e-8 ute=-2.093499336e+00 lute=1.575544871e-07 wute=1.182086919e-05 pute=-4.259368433e-12 ua1=-3.367642224e-10 lua1=3.417072675e-16 wua1=2.454381866e-14 pua1=-8.711290378e-21 ub1=-1.075982408e-19 lub1=-1.809441990e-25 wub1=-1.121342091e-23 pub1=2.837218933e-30 uc1=1.802069720e-11 luc1=9.801780433e-18 wuc1=6.970910250e-16 puc1=-4.749569907e-22 kt1l=0.0 prt=0.0 tvoff=1.074871566e-03 ltvoff=-2.562295865e-10 wtvoff=-4.271056080e-09 ptvoff=3.609895022e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.6 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.547564871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.310308032e-09 wvth0=4.581457956e-07 pvth0=-1.310578374e-13 k1=5.706865460e-01 lk1=-7.045806481e-09 wk1=-2.080563774e-06 pk1=7.047260171e-13 k2=-4.668578416e-02 lk2=1.681842852e-09 wk2=6.010738037e-07 pk2=-1.682189850e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.591628369e-01 ldsub=-4.146408340e-09 wdsub=8.373358603e-08 pdsub=4.147263827e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.608891738e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.663651286e-10 wvoff=-3.589206583e-07 pvoff=9.665645090e-14 nfactor=2.820951068e+00 lnfactor=-5.983427045e-09 wnfactor=-1.685454455e-06 pnfactor=5.984661546e-13 eta0=-3.645268133e-02 weta0=3.696030541e-6 etab=-5.482800931e-04 letab=1.473784182e-11 wetab=4.759884163e-09 petab=-1.474088253e-15 u0=3.111783475e-02 lu0=1.264910037e-10 wu0=-3.122991688e-08 pu0=-1.265171014e-14 ua=-9.035873898e-10 lua=1.328153242e-17 wua=-2.102231667e-15 pua=-1.328427266e-21 ub=1.847142908e-18 lub=-8.988261670e-27 wub=1.092934622e-24 pub=8.990116128e-31 uc=7.378357019e-11 luc=-4.694495689e-20 wuc=5.305392466e-17 puc=4.695464258e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.851921306e+04 lvsat=-3.172166976e-04 wvsat=1.481092453e-01 pvsat=3.172821457e-8 a0=1.075417795e+00 wa0=2.980835418e-6 ags=5.802298781e-01 lags=3.141072004e-08 wags=1.131894703e-05 pags=-3.141720070e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.213177679e-03 lketa=2.988377852e-10 wketa=-1.340774250e-07 pketa=-2.988994414e-14 dwg=0.0 dwb=0.0 pclm=5.536471621e-01 lpclm=3.180973941e-09 wpclm=5.503973278e-07 ppclm=-3.181630240e-13 pdiblc1=2.929611003e-01 lpdiblc1=2.251119149e-08 wpdiblc1=9.705892081e-06 ppdiblc1=-2.251583600e-12 pdiblc2=4.866013531e-03 lpdiblc2=2.260401717e-11 wpdiblc2=-5.353117278e-09 ppdiblc2=-2.260868083e-15 pdiblcb=-3.656432464e-02 lpdiblcb=5.105487427e-09 wpdiblcb=1.156671059e-06 ppdiblcb=-5.106540791e-13 drout=5.936065733e-01 ldrout=-1.279556685e-08 wdrout=-3.361350705e-06 pdrout=1.279820683e-12 pscbe1=8.318856122e+08 lpscbe1=-6.105648330e+00 wpscbe1=-3.189219080e+03 ppscbe1=6.106908047e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.149599339e-07 lalpha0=8.577218877e-14 walpha0=6.450930020e-11 palpha0=-8.578988529e-18 alpha1=0.85 beta0=1.350598378e+01 lbeta0=-8.347471943e-09 wbeta0=3.540892632e-05 pbeta0=8.349194194e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.284076625e-01 lkt1=3.806661637e-10 wkt1=4.428576060e-07 pkt1=-3.807447027e-14 kt2=-4.745543019e-02 lkt2=9.887424799e-11 wkt2=1.007052923e-07 pkt2=-9.889464773e-15 at=1.179932801e+05 lat=7.020959860e-04 wat=-3.053910028e-01 pat=-7.022408425e-8 ute=-1.704349548e+00 lute=-1.424969596e-08 wute=-1.055262843e-06 pute=1.425263595e-12 ua1=4.567635353e-10 lua1=-8.624128096e-18 wua1=2.858236063e-15 pua1=8.625907426e-22 ub1=-4.924731976e-19 lub1=-1.102729379e-26 wub1=-7.285183007e-24 pub1=1.102956894e-30 uc1=4.622357190e-11 luc1=-2.649393909e-18 wuc1=-9.789554269e-16 puc1=2.649940532e-22 kt1l=0.0 prt=0.0 tvoff=4.466454610e-04 ltvoff=2.112344368e-11 wtvoff=8.691246708e-09 ptvoff=-2.112780187e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.7 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.510514691e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.019767105e-09 wvth0=8.287240357e-07 pvth0=-2.020183823e-13 k1=5.502646663e-01 lk1=-3.135302414e-09 wk1=-3.795445444e-08 pk1=3.135949290e-13 k2=-4.045406726e-02 lk2=4.885563109e-10 wk2=-2.222645860e-08 pk2=-4.886571099e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.166789622e-01 ldsub=3.988658889e-09 wdsub=4.332997582e-06 pdsub=-3.989481829e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.703927872e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.534437798e-10 wvoff=5.916367565e-07 pvoff=-8.536198623e-14 nfactor=2.742020436e+00 lnfactor=9.130683879e-09 wnfactor=6.209237203e-06 pnfactor=-9.132567721e-13 eta0=-9.659088373e-02 leta0=1.151562382e-08 weta0=9.711091552e-06 peta0=-1.151799973e-12 etab=-4.069996608e-03 letab=6.890972504e-10 wetab=3.570041957e-07 petab=-6.892394249e-14 u0=3.284197820e-02 lu0=-2.036583298e-10 wu0=-2.036798349e-07 pu0=2.037003486e-14 ua=-6.476465638e-10 lua=-3.572755258e-17 wua=-2.770159483e-14 pua=3.573492389e-21 ub=1.649677481e-18 lub=2.882360319e-26 wub=2.084355148e-23 pub=-2.882955007e-30 uc=7.377567729e-11 luc=-4.543357708e-20 wuc=5.384337749e-17 puc=4.544295093e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.793719399e+04 lvsat=-2.057681939e-04 wvsat=2.063231605e-01 pvsat=2.058106480e-8 a0=1.075417795e+00 wa0=2.980835418e-6 ags=9.054765746e-01 lags=-3.086946889e-08 wags=-2.121243311e-05 pags=3.087583787e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.683864836e-03 lketa=1.722178429e-11 wketa=-2.811764840e-07 pketa=-1.722533749e-15 dwg=0.0 dwb=0.0 pclm=5.538089467e-01 lpclm=3.149994444e-09 wpclm=5.342155237e-07 ppclm=-3.150644351e-13 pdiblc1=4.441554486e-01 lpdiblc1=-6.440409498e-09 wpdiblc1=-5.416662196e-06 ppdiblc1=6.441738284e-13 pdiblc2=5.808102089e-03 lpdiblc2=-1.577927525e-10 wpdiblc2=-9.958141025e-08 ppdiblc2=1.578253083e-14 pdiblcb=8.262579618e-03 lpdiblcb=-3.478237161e-09 wpdiblcb=-3.326944235e-06 ppdiblcb=3.478954791e-13 drout=4.896939158e-01 ldrout=7.102252282e-09 wdrout=7.032058972e-06 pdrout=-7.103717619e-13 pscbe1=7.994623781e+08 lpscbe1=1.029470667e-01 wpscbe1=5.377328201e+01 ppscbe1=-1.029683068e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.116263740e-07 lalpha0=6.598525873e-14 walpha0=5.417381224e-11 palpha0=-6.599887281e-18 alpha1=8.946892610e-01 lalpha1=-8.557367830e-09 walpha1=-4.469848128e-06 palpha1=8.559133387e-13 beta0=1.292169122e+01 lbeta0=1.035363736e-07 wbeta0=9.385023765e-05 pbeta0=-1.035577352e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.221573236e-01 lkt1=-8.161862395e-10 wkt1=-1.823052455e-07 pkt1=8.163546351e-14 kt2=-4.644251018e-02 lkt2=-9.508575335e-11 wkt2=-6.076073935e-10 pkt2=9.510537145e-15 at=1.229755015e+05 lat=-2.519296616e-04 wat=-8.037159363e-01 pat=2.519816397e-8 ute=-1.903959091e+00 lute=2.397273693e-08 wute=1.890980977e-05 pute=-2.397768299e-12 ua1=1.476705289e-10 lua1=5.056285533e-17 wua1=3.377391391e-14 pua1=-5.057328745e-21 ub1=-3.293871992e-19 lub1=-4.225597929e-26 wub1=-2.359714764e-23 pub1=4.226469754e-30 uc1=3.783361613e-11 luc1=-1.042834837e-18 wuc1=-1.397867478e-16 puc1=1.043049995e-22 kt1l=0.0 prt=0.0 tvoff=6.618992138e-04 ltvoff=-2.009463643e-11 wtvoff=-1.283856969e-08 ptvoff=2.009878235e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.8 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.473610650e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.468099541e-09 wvth0=1.197840589e-06 pvth0=-2.468608759e-13 k1=5.281406079e-01 lk1=-4.475390587e-10 wk1=2.174907846e-06 pk1=4.476313949e-14 k2=-3.013986029e-02 lk2=-7.644754372e-10 wk2=-1.053859958e-06 pk2=7.646331638e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.328412677e-01 ldsub=2.025165043e-09 wdsub=2.716433572e-06 pdsub=-2.025582875e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=4.156859372e-03 lcdscd=1.510242328e-10 wcdscd=1.243397528e-07 pcdscd=-1.510553921e-14 cit=0.0 voff='-2.659283894e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.110819521e-10 wvoff=1.451048699e-07 pvoff=-3.111461346e-14 nfactor=2.811345204e+00 lnfactor=7.086951962e-10 wnfactor=-7.246698378e-07 pnfactor=-7.088414142e-14 eta0=-8.753769020e-03 leta0=8.446441062e-10 weta0=9.255678258e-07 peta0=-8.448183732e-14 etab=-1.673778762e-03 letab=3.979903292e-10 wetab=1.173329724e-07 petab=-3.980724426e-14 u0=2.849673133e-02 lu0=3.242283319e-10 wu0=2.309345037e-07 pu0=-3.242952267e-14 ua=-1.327109946e-09 lua=4.681773591e-17 wua=4.025876211e-14 pua=-4.682739535e-21 ub=2.219978211e-18 lub=-4.045995132e-26 wub=-3.619828798e-23 pub=4.046829902e-30 uc=6.574233499e-11 luc=9.305050463e-19 wuc=8.573433520e-16 puc=-9.306970281e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.706851076e+04 lvsat=-1.002353427e-04 wvsat=2.932094065e-01 pvsat=1.002560232e-8 a0=1.075417795e+00 wa0=2.980835418e-6 ags=6.513775930e-01 wags=4.202707627e-6 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.704117229e-02 lketa=-1.726990070e-09 wketa=-1.717203450e-06 pketa=1.727346382e-13 dwg=0.0 dwb=0.0 pclm=5.528169047e-01 lpclm=3.270513664e-09 wpclm=6.334401962e-07 ppclm=-3.271188436e-13 pdiblc1=3.938665019e-01 lpdiblc1=-3.310065232e-10 wpdiblc1=-3.867299674e-07 ppdiblc1=3.310748165e-14 pdiblc2=4.675550531e-03 lpdiblc2=-2.020359396e-11 wpdiblc2=1.369711228e-08 ppdiblc2=2.020776237e-15 pdiblcb=-4.902386720e-04 lpdiblcb=-2.414892278e-09 wpdiblcb=-2.451481818e-06 ppdiblcb=2.415390519e-13 drout=5.066442075e-01 ldrout=5.043029150e-09 wdrout=5.336680087e-06 pdrout=-5.044069627e-13 pscbe1=7.990756346e+08 lpscbe1=1.499309852e-01 wpscbe1=9.245560931e+01 ppscbe1=-1.499619189e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.617456841e-08 lalpha0=-5.648865656e-16 walpha0=-6.175842348e-13 palpha0=5.650031130e-20 alpha1=7.457250577e-01 lalpha1=9.539697373e-09 walpha1=1.042964563e-05 palpha1=-9.541665603e-13 beta0=1.351149975e+01 lbeta0=3.188289359e-08 wbeta0=3.485721495e-05 pbeta0=-3.188947167e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.188134799e-01 lkt1=-1.222416430e-09 wkt1=-5.167586012e-07 pkt1=1.222668639e-13 kt2=-4.567643327e-02 lkt2=-1.881533726e-10 wkt2=-7.723110393e-08 pkt2=1.881921924e-14 at=1.201564742e+05 lat=9.054269131e-05 wat=-5.217550423e-01 pat=-9.056137208e-9 ute=-1.286620494e+00 lute=-5.102525985e-08 wute=-4.283678685e-05 pute=5.103578738e-12 ua1=1.148833628e-09 lua1=-7.106444492e-17 wua1=-6.636305199e-14 pua1=7.107910694e-21 ub1=-1.012443069e-18 lub1=4.072574614e-26 wub1=4.472253217e-23 pub1=-4.073414867e-30 uc1=3.550642909e-11 luc1=-7.601141930e-19 wuc1=9.297997050e-17 puc1=7.602710198e-23 kt1l=0.0 prt=0.0 tvoff=2.587882778e-04 ltvoff=2.887769874e-11 wtvoff=2.748084090e-08 ptvoff=-2.888365679e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.9 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.413635332e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.749623453e-08 wvth0=-6.848859382e-09 pvth0=6.844851840e-13 k1=5.418278423e-01 lk1=-9.616293131e-08 wk1=-6.755198265e-09 pk1=6.751245528e-13 k2=-3.150321751e-02 lk2=1.948924088e-08 wk2=1.369068979e-09 pk2=-1.368267882e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.553056256e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.639672501e-07 wvoff=-3.961724686e-08 pvoff=3.959406523e-12 nfactor=3.418446533e+00 lnfactor=-7.368251346e-05 wnfactor=-5.176006807e-06 pnfactor=5.172978119e-10 eta0=0.08 etab=-0.07 u0=3.205529497e-02 lu0=5.408883467e-08 wu0=3.799601334e-09 pu0=-3.797378035e-13 ua=-7.341927684e-10 lua=-2.379836807e-15 wua=-1.671774066e-16 pua=1.670795844e-20 ub=1.661783026e-18 lub=7.367863613e-24 wub=5.175734434e-25 pub=-5.172705905e-29 uc=4.770329823e-11 luc=1.537801416e-16 wuc=1.080265890e-17 puc=-1.079633783e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.279687104e+00 la0=-1.455251685e-07 wa0=-1.022276830e-08 pa0=1.021678655e-12 ags=4.491558820e-01 lags=6.202486556e-07 wags=4.357087065e-08 pags=-4.354537560e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=7.886878719e-25 lb1=1.317882931e-28 wb1=9.257788177e-30 pb1=-9.252371074e-34 keta=-7.162882048e-03 lketa=-1.630763169e-07 wketa=-1.145569127e-08 pketa=1.144898809e-12 dwg=0.0 dwb=0.0 pclm=5.795731508e-02 lpclm=-3.162280048e-06 wpclm=-2.221420292e-07 ppclm=2.220120450e-11 pdiblc1=0.39 pdiblc2=3.148691893e-03 lpdiblc2=-7.518917112e-09 wpdiblc2=-5.281845627e-10 ppdiblc2=5.278755008e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.170395671e+08 lpscbe1=3.761257139e+03 wpscbe1=2.642186272e+02 ppscbe1=-2.640640223e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.201446967e-01 lkt1=7.110533590e-07 wkt1=4.994966721e-08 pkt1=-4.992043966e-12 kt2=-4.543608648e-02 lkt2=1.226776545e-08 wkt2=8.617789285e-10 pkt2=-8.612746672e-14 at=140000.0 ute=-1.857389725e+00 lute=4.396398517e-06 wute=3.088356732e-07 pute=-3.086549611e-11 ua1=3.028581411e-10 lua1=7.311904902e-15 wua1=5.136424881e-16 pua1=-5.133419353e-20 ub1=-5.509084302e-19 lub1=-8.865966113e-24 wub1=-6.228112858e-25 pub1=6.224468540e-29 uc1=1.657886115e-11 luc1=-7.487097943e-17 wuc1=-5.259493481e-18 puc1=5.256415941e-22 kt1l=0.0 prt=0.0 tvoff=1.497522209e-03 ltvoff=-5.279930782e-08 wtvoff=-3.709015394e-09 ptvoff=3.706845101e-13 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.10 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.364744174e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.747582355e-8 k1=5.370055873e-01 wk1=2.710007976e-8 k2=-3.052589612e-02 wk2=-5.492344868e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.835867301e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=1.589339806e-7 nfactor=-2.764894144e-01 wnfactor=2.076477874e-5 eta0=0.08 etab=-0.07 u0=3.476767231e-02 wu0=-1.524300179e-8 ua=-8.535337647e-10 wua=6.706718110e-16 ub=2.031257177e-18 wub=-2.076368605e-24 uc=5.541486704e-11 wuc=-4.333742790e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.272389495e+00 wa0=4.101105926e-8 ags=4.802593141e-01 wags=-1.747948800e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=7.397437744e-24 wb1=-3.713981266e-29 keta=-1.534062351e-02 wketa=4.595722212e-8 dwg=0.0 dwb=0.0 pclm=-1.006206389e-01 wpclm=8.911754287e-7 pdiblc1=0.39 pdiblc2=2.771642905e-03 wpdiblc2=2.118937627e-9 pdiblcb=-0.025 drout=0.56 pscbe1=9.056542541e+08 wpscbe1=-1.059975680e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.844877071e-01 wkt1=-2.003849350e-7 kt2=-4.482089835e-02 wkt2=-3.457230533e-9 at=140000.0 ute=-1.636924785e+00 wute=-1.238967540e-6 ua1=6.695261467e-10 wua1=-2.060598646e-15 ub1=-9.955074993e-19 wub1=2.498555166e-24 uc1=1.282432754e-11 wuc1=2.109970533e-17 kt1l=0.0 prt=0.0 tvoff=-1.150189592e-03 wtvoff=1.487959481e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.11 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.219179249e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.156001811e-07 wvth0=6.887682548e-08 pvth0=-3.287854772e-13 k1=5.247275001e-01 lk1=9.750625747e-08 wk1=5.001754881e-08 pk1=-1.819987596e-13 k2=-2.098959161e-02 lk2=-7.573242878e-08 wk2=-1.913369715e-08 pk2=1.083326081e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.896740758e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.834257061e-08 wvoff=2.233272999e-07 pvoff=-5.113786434e-13 nfactor=-2.661313226e+00 lnfactor=1.893904491e-05 wnfactor=3.747800200e-05 pnfactor=-1.327278286e-10 eta0=0.08 etab=-0.07 u0=3.642278220e-02 lu0=-1.314403201e-08 wu0=-2.675105629e-08 pu0=9.139105377e-14 ua=-8.963917912e-10 lua=3.403564175e-16 wua=9.352766592e-16 pua=-2.101355698e-21 ub=2.240454184e-18 lub=-1.661335101e-24 wub=-3.613967779e-24 pub=1.221082231e-29 uc=1.759490555e-10 luc=-9.572205699e-16 wuc=-8.456555022e-16 puc=6.371597755e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.694078634e+00 la0=-3.348838398e-06 wa0=-2.170833996e-06 pa0=1.756533654e-11 ags=6.127202719e-01 lags=-1.051936842e-06 wags=-1.199038996e-06 pags=8.134020310e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=1.468666207e-23 lb1=-5.788727294e-29 wb1=-7.373632556e-29 pb1=2.906306949e-34 keta=-2.855092721e-02 lketa=1.049094419e-07 wketa=9.157211667e-08 pketa=-3.622500464e-13 dwg=0.0 dwb=0.0 pclm=-1.017522331e+00 lpclm=7.281561951e-06 wpclm=3.449493382e-06 ppclm=-2.031684621e-11 pdiblc1=0.39 pdiblc2=2.811135398e-03 lpdiblc2=-3.136290773e-10 wpdiblc2=1.723189895e-09 ppdiblc2=3.142825071e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.007119366e+09 lpscbe1=-8.057837632e+02 wpscbe1=-2.085885908e+03 ppscbe1=8.147251718e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.592309989e-01 lkt1=-2.005757943e-07 wkt1=-3.631061549e-07 pkt1=1.292248289e-12 kt2=-3.210563747e-02 lkt2=-1.009780663e-07 wkt2=-8.496849217e-08 pkt2=6.473205431e-13 at=140000.0 ute=-1.115603560e+00 lute=-4.140065214e-06 wute=-4.623638378e-06 pute=2.687931607e-11 ua1=1.925939265e-09 lua1=-9.977787188e-15 wua1=-9.518857161e-15 pua1=5.922965558e-20 ub1=-2.199445576e-18 lub1=9.561057381e-24 wub1=9.167172927e-24 pub1=-5.295873459e-29 uc1=-2.776324147e-11 luc1=3.223256111e-16 wuc1=2.055484280e-16 puc1=-1.464796949e-21 kt1l=0.0 prt=0.0 tvoff=-2.894179300e-03 ltvoff=1.384986984e-08 wtvoff=2.830557157e-08 ptvoff=-1.066222065e-13 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.12 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.439420063e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.879257239e-08 wvth0=-3.250360229e-08 pvth0=7.080405949e-14 k1=5.754007465e-01 lk1=-1.022216339e-07 wk1=-1.773635804e-07 pk1=7.142207778e-13 k2=-5.285786008e-02 lk2=4.987590525e-08 wk2=1.085186711e-07 pk2=-3.948074142e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.287789319e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.916747864e-07 wvoff=-2.451127946e-07 pvoff=1.334971431e-12 nfactor=2.695058914e+00 lnfactor=-2.173020889e-06 wnfactor=-8.755341785e-07 pnfactor=1.844209736e-11 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374642839e-01 letab=2.659095304e-07 wetab=-1.182120578e-11 petab=4.659311709e-17 u0=3.545030617e-02 lu0=-9.311031345e-09 wu0=-8.053854486e-09 pu0=1.769629460e-14 ua=-4.143713417e-10 lua=-1.559520436e-15 wua=-1.204535523e-15 pua=6.332684062e-21 ub=1.399856672e-18 lub=1.651868223e-24 wub=1.658959981e-24 pub=-8.572348631e-30 uc=-2.100382789e-10 luc=5.641431046e-16 wuc=1.561623780e-15 puc=-3.116659834e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=4.925112385e-01 la0=1.387122670e-06 wa0=5.198000524e-06 pa0=-1.147882156e-11 ags=-7.062784917e-02 lags=1.641470210e-06 wags=2.259093814e-06 pags=-5.496161747e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.682948282e-07 lketa=-7.621792194e-09 wketa=-2.655029092e-08 pketa=1.033277694e-13 dwg=0.0 dwb=0.0 pclm=8.375014444e-01 lpclm=-2.998828922e-08 wpclm=-1.568597601e-06 ppclm=-5.381108521e-13 pdiblc1=0.39 pdiblc2=1.353724391e-03 lpdiblc2=5.430736003e-09 wpdiblc2=4.586723084e-10 ppdiblc2=8.126903435e-15 pdiblcb=-0.025 drout=0.56 pscbe1=8.052871584e+08 lpscbe1=-1.026494406e+01 wpscbe1=-3.711919361e+01 ppscbe1=7.206639473e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.047546705e-01 lkt1=-2.114488008e-08 wkt1=-1.266494896e-08 pkt1=-8.901081765e-14 kt2=-5.828982076e-02 lkt2=2.226525553e-09 wkt2=8.332428097e-08 pkt2=-1.600306609e-14 at=1.673241718e+05 lat=-1.076978404e-01 wat=-2.104330658e-02 pat=8.294189826e-8 ute=-2.534178812e+00 lute=1.451229284e-06 wute=3.838355419e-06 pute=-6.473514011e-12 ua1=-1.722329642e-09 lua1=4.401813633e-15 wua1=1.126158851e-14 pua1=-2.267618012e-20 ub1=1.240467215e-18 lub1=-3.997310726e-24 wub1=-1.013826331e-23 pub1=2.313337205e-29 uc1=6.758595409e-11 luc1=-5.349190836e-17 wuc1=-3.027950207e-16 puc1=5.388316375e-22 kt1l=0.0 prt=0.0 tvoff=7.623177698e-04 ltvoff=-5.621621641e-10 wtvoff=2.057709918e-09 ptvoff=-3.166627270e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.13 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.420624745e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.244165713e-08 wvth0=2.748728890e-08 pvth0=-4.566741589e-14 k1=4.361991255e-01 lk1=1.680363645e-07 wk1=5.750620115e-07 pk1=-7.466029749e-13 k2=8.295027818e-03 lk2=-6.885157047e-08 wk2=-2.787552946e-07 pk2=3.570795683e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.113048857e+00 ldsub=-1.656182414e-06 wdsub=-5.988942104e-06 pdsub=1.162744725e-11 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.808720934e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.036119574e-07 wvoff=8.760463320e-07 pvoff=-8.417433173e-13 nfactor=-1.859309060e-01 lnfactor=3.420380513e-06 wnfactor=2.077930357e-05 pnfactor=-2.360046695e-11 eta0=-6.227434766e-03 leta0=1.306122041e-08 weta0=3.380463323e-08 peta0=-6.563122215e-14 etab=-9.503404713e-04 letab=8.696204559e-10 wetab=1.912912609e-09 petab=-3.690250638e-15 u0=3.467445811e-02 lu0=-7.804733206e-09 wu0=4.159495940e-09 pu0=-6.015754263e-15 ua=-9.507846956e-10 lua=-5.180814192e-16 wua=3.595714803e-15 pua=-2.986934743e-21 ub=2.144869552e-18 lub=2.054361479e-25 wub=-4.851760495e-24 pub=4.068124022e-30 uc=7.465980580e-11 luc=1.140575896e-17 wuc=8.641490596e-17 puc=-2.525624581e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.205199566e+04 lvsat=1.125052391e-01 wvsat=2.726521308e-01 pvsat=-5.293502948e-7 a0=2.337983204e+00 la0=-2.195835314e-06 wa0=-8.025894747e-06 pa0=1.419518598e-11 ags=1.467233020e+00 lags=-1.344265137e-06 wags=-7.211998617e-06 pags=1.289183161e-11 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.933150141e-02 lketa=-1.033991207e-07 wketa=8.203966215e-08 pketa=-1.074981043e-13 dwg=0.0 dwb=0.0 pclm=1.091728878e+00 lpclm=-5.235672927e-07 wpclm=-2.632092630e-06 ppclm=1.526649858e-12 pdiblc1=-1.712753477e-01 lpdiblc1=1.089708230e-06 wpdiblc1=1.844118494e-06 ppdiblc1=-3.580330238e-12 pdiblc2=6.735720638e-03 lpdiblc2=-5.018334363e-09 wpdiblc2=-8.207294483e-09 ppdiblc2=2.495175664e-14 pdiblcb=-4.813289512e-02 lpdiblcb=4.491219201e-08 wpdiblcb=-1.571733722e-09 ppdiblcb=3.051499017e-15 drout=8.424458000e-01 ldrout=-5.483645665e-7 pscbe1=2.285248550e+09 lpscbe1=-2.883589266e+03 wpscbe1=-6.865179715e+03 ppscbe1=1.332865030e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=4.088343835e-07 lalpha0=-7.355016519e-13 walpha0=-1.991130458e-11 palpha0=3.865751909e-17 alpha1=8.179894760e-01 lalpha1=6.214798420e-8 beta0=1.190487019e+01 lbeta0=3.795857156e-06 wbeta0=-4.596192808e-06 pbeta0=8.923443991e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.581993095e-01 lkt1=8.261713836e-08 wkt1=-9.877683398e-08 pkt1=7.817420155e-14 kt2=-8.619110695e-02 lkt2=5.639648208e-08 wkt2=1.464126456e-07 pkt2=-1.384882427e-13 at=1.545264453e+05 lat=-8.285123375e-02 wat=6.297333936e-02 pat=-8.017524359e-8 ute=-2.534936483e+00 lute=1.452700291e-06 wute=2.837038937e-07 pute=4.277921599e-13 ua1=-8.022069977e-10 lua1=2.615408400e-15 wua1=-2.322012134e-15 pua1=3.696190366e-21 ub1=-3.714809550e-19 lub1=-8.677359211e-25 wub1=4.604204679e-24 pub1=-5.488923150e-30 uc1=1.270684976e-11 luc1=5.305510440e-17 wuc1=3.815695325e-17 puc1=-1.231218466e-22 kt1l=0.0 prt=0.0 tvoff=-2.239112263e-04 ltvoff=1.352587625e-09 wtvoff=3.949816576e-09 ptvoff=-6.840125857e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.14 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.822414253e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.386262557e-09 wvth0=-1.056398641e-07 pvth0=7.966993488e-14 k1=7.104378696e-01 lk1=-9.015557370e-08 wk1=-2.833974873e-07 pk1=6.162462481e-14 k2=-1.085580177e-01 lk2=4.116393599e-08 wk2=1.658085416e-07 pk2=-6.147105955e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.652016335e+00 ldsub=9.470877538e-07 wdsub=1.258358629e-05 pdsub=-5.858328221e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.157208325e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.187564275e-08 wvoff=-3.451430200e-07 pvoff=3.079893610e-13 nfactor=5.718571529e+00 lnfactor=-2.138625867e-06 wnfactor=-1.976539436e-05 pnfactor=1.457179852e-11 eta0=-4.182599245e-01 leta0=4.009840410e-07 weta0=-6.760926646e-08 peta0=2.984854461e-14 etab=2.257051638e-04 letab=-2.376100449e-10 wetab=-3.778540395e-09 petab=1.668172685e-15 u0=3.034164638e-02 lu0=-3.725451627e-09 wu0=-1.021848342e-08 pu0=7.520912013e-15 ua=-1.291682198e-09 lua=-1.971311930e-16 wua=-5.044163920e-17 pua=4.458705014e-22 ub=2.336274434e-18 lub=2.523113104e-26 wub=-2.499146522e-25 pub=-2.644494133e-31 uc=8.763791370e-11 luc=-8.129479379e-19 wuc=-3.235164034e-16 puc=1.333821307e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.854494372e+05 lvsat=-4.133116447e-02 wvsat=-6.525619196e-01 pvsat=3.417257807e-7 a0=-1.313771719e+00 la0=1.242240821e-06 wa0=1.327783687e-05 pa0=-5.861979088e-12 ags=-1.029486580e+00 lags=1.006361412e-06 wags=1.220367177e-05 pags=-5.387750233e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-7.935737222e-02 lketa=1.775965215e-08 wketa=-1.366379865e-07 pketa=9.838384046e-14 dwg=0.0 dwb=0.0 pclm=2.848871364e-01 lpclm=2.360629113e-07 wpclm=-1.486087973e-07 ppclm=-8.115154019e-13 pdiblc1=7.045990381e-01 lpdiblc1=2.650847577e-07 wpdiblc1=-1.797308830e-06 ppdiblc1=-1.519773930e-13 pdiblc2=-1.316612295e-03 lpdiblc2=2.562824361e-09 wpdiblc2=4.103947058e-08 ppdiblc2=-2.141338322e-14 pdiblcb=2.126579023e-02 lpdiblcb=-2.042569867e-08 wpdiblcb=3.143467444e-09 ppdiblcb=-1.387796868e-15 drout=9.768540291e-01 ldrout=-6.749080325e-07 wdrout=-6.512799530e-06 pdrout=6.131709578e-12 pscbe1=-1.429156617e+09 lpscbe1=6.134711971e+02 wpscbe1=1.000836168e+04 ppscbe1=-2.557552689e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.923174788e-05 lalpha0=1.775583158e-11 walpha0=1.327247809e-10 palpha0=-1.050472185e-16 alpha1=9.140210480e-01 lalpha1=-2.826439640e-08 walpha1=3.552713679e-21 beta0=2.458676570e+00 lbeta0=1.268931620e-05 wbeta0=8.606620946e-05 pbeta0=-7.643393847e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.687837559e-01 lkt1=-1.566353585e-09 wkt1=-2.256275305e-09 pkt1=-1.269855316e-14 kt2=-1.821576988e-02 lkt2=-7.601346121e-09 wkt2=2.709858025e-09 pkt2=-3.194080083e-15 at=7.900862825e+04 lat=-1.175226621e-02 wat=-4.821526100e-02 pat=2.450726701e-8 ute=-7.067122344e-01 lute=-2.685472438e-07 wute=2.084747293e-06 pute=-1.267864986e-12 ua1=2.530268617e-09 lua1=-5.220707360e-16 wua1=4.415436167e-15 pua1=-2.647022885e-21 ub1=-1.237565052e-18 lub1=-5.232986928e-26 wub1=-3.280339758e-24 pub1=1.934265054e-30 uc1=1.442870135e-10 luc1=-7.082577767e-17 wuc1=-1.893783160e-16 puc1=9.109942387e-23 kt1l=0.0 prt=0.0 tvoff=2.270495240e-03 ltvoff=-9.958611414e-10 wtvoff=-1.266508990e-08 ptvoff=8.802575984e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.15 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.016963394e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.397533475e-08 wvth0=1.285983665e-07 pvth0=-2.374296458e-14 k1=3.171094464e-01 lk1=8.349341856e-08 wk1=-3.002922739e-07 pk1=6.908343654e-14 k2=2.780929504e-02 lk2=-1.904032346e-08 wk2=7.807126687e-08 pk2=-2.273628109e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.050777091e-01 ldsub=3.890953274e-08 wdsub=-9.406810354e-07 pdsub=1.124464649e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.461848609e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.987099931e-08 wvoff=9.419721720e-07 pvoff=-2.602539767e-13 nfactor=-1.450591710e+00 lnfactor=1.026459335e-06 wnfactor=2.830347546e-05 pnfactor=-6.649934537e-12 eta0=0.49 etab=-2.706292950e-04 letab=-1.848533005e-11 wetab=2.810600086e-09 petab=-1.240840589e-15 u0=2.418140125e-02 lu0=-1.005789641e-09 wu0=1.746823013e-08 pu0=-4.702384407e-15 ua=-1.411309201e-09 lua=-1.443175461e-16 wua=1.462296327e-15 pua=-2.219821323e-22 ub=2.102599493e-18 lub=1.283953463e-25 wub=-7.005320487e-25 pub=-6.550814140e-32 uc=1.571267704e-11 luc=3.094103709e-17 wuc=4.607482954e-16 puc=-2.128597541e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.260003180e+04 lvsat=1.290512811e-02 wvsat=2.598719587e-01 pvsat=-6.110100252e-8 a0=1.5 ags=2.192470828e+00 lags=-4.160876762e-07 wags=-3.374750193e-12 pags=1.489904963e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.761266914e-02 lketa=-5.084909831e-09 wketa=6.829823754e-08 pketa=7.907366649e-15 dwg=0.0 dwb=0.0 pclm=1.157511655e+00 lpclm=-1.491885967e-07 wpclm=-3.689113052e-06 ppclm=7.515676594e-13 pdiblc1=2.947449378e+00 lpdiblc1=-7.251022676e-07 wpdiblc1=-8.930293268e-06 ppdiblc1=2.997135375e-12 pdiblc2=5.965945468e-03 lpdiblc2=-6.523229356e-10 wpdiblc2=-1.307533463e-08 ppdiblc2=2.477545680e-15 pdiblcb=5.127410957e-01 lpdiblcb=-2.374051654e-07 wpdiblcb=-2.699800153e-06 ppdiblcb=1.191923970e-12 drout=-1.740506618e+00 ldrout=5.247686503e-07 wdrout=1.302559906e-05 pdrout=-2.494219862e-12 pscbe1=-6.826809653e+08 lpscbe1=2.839126473e+02 wpscbe1=7.443995500e+03 ppscbe1=-1.425420922e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.861538074e-05 lalpha0=-7.782865843e-12 walpha0=-2.109124849e-10 palpha0=4.666382343e-17 alpha1=0.85 beta0=4.098154398e+01 lbeta0=-4.317990442e-06 wbeta0=-1.574868709e-04 pbeta0=3.109133676e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.227247028e-01 lkt1=-2.190078067e-08 wkt1=-2.991035628e-07 pkt1=1.183553684e-13 kt2=-5.987419801e-03 lkt2=-1.299999148e-08 wkt2=-1.904263484e-07 pkt2=8.207285114e-14 at=7.508357758e+04 lat=-1.001941130e-02 wat=-4.137772372e-03 pat=5.047672862e-9 ute=-1.220298243e+00 lute=-4.180621117e-08 wute=-4.453608926e-06 pute=1.618727748e-12 ua1=1.695712953e-09 lua1=-1.536260941e-16 wua1=-5.839971865e-15 pua1=1.880596185e-21 ub1=-1.994757491e-18 lub1=2.819599921e-25 wub1=3.261802178e-24 pub1=-9.539990204e-31 uc1=-1.178169179e-10 luc1=4.488943860e-17 wuc1=1.727124851e-16 puc1=-6.875859554e-23 kt1l=0.0 prt=0.0 tvoff=1.916901178e-04 ltvoff=-7.809778338e-11 wtvoff=1.048119435e-08 ptvoff=-1.416184465e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.16 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.567769459e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.452249976e-08 wvth0=8.646437025e-08 pvth0=-1.567489418e-14 k1=5.233086898e-01 lk1=4.400915023e-08 wk1=1.512935363e-07 pk1=-1.738892391e-14 k2=-3.862583202e-02 lk2=-6.318926721e-09 wk2=-3.506182542e-08 pk2=-1.072877775e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=9.554854829e-01 ldsub=-6.648585023e-08 wdsub=-8.538911190e-07 pdsub=9.582741101e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='8.459525931e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.176596279e-08 wvoff=-1.900603682e-06 pvoff=2.840595034e-13 nfactor=5.457562658e+00 lnfactor=-2.963555124e-07 wnfactor=-1.285558541e-05 pnfactor=1.231449393e-12 eta0=1.315407875e+00 leta0=-1.580540523e-07 weta0=-2.020321159e-07 peta0=3.868632174e-14 etab=6.198423664e-02 letab=-1.193942059e-08 wetab=-1.067382680e-07 petab=1.973623396e-14 u0=4.544915689e-03 lu0=2.754322432e-09 wu0=-5.016572301e-09 pu0=-3.968595279e-16 ua=-4.589156849e-09 lua=4.641957886e-16 wua=-2.970159713e-17 pua=6.371458218e-23 ub=4.322530794e-18 lub=-2.966904188e-25 wub=2.078431984e-24 pub=-5.976408481e-31 uc=3.130273050e-10 luc=-2.599055176e-17 wuc=-1.625854256e-15 puc=1.866954221e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.705514603e+04 lvsat=1.013717611e-02 wvsat=2.125156947e-01 pvsat=-5.203294095e-8 a0=1.5 ags=-2.115967244e+00 lags=4.089178967e-07 wags=1.205267926e-11 pags=-1.464231792e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.008928720e-01 lketa=8.947223101e-09 wketa=4.459976694e-07 pketa=-6.441678675e-14 dwg=0.0 dwb=0.0 pclm=1.003620026e+00 lpclm=-1.197205044e-07 wpclm=-2.623742536e-06 ppclm=5.475641208e-13 pdiblc1=-2.944097377e+00 lpdiblc1=4.030464544e-07 wpdiblc1=1.837101401e-05 ppdiblc1=-2.230682752e-12 pdiblc2=-6.305032684e-03 lpdiblc2=1.697397587e-09 wpdiblc2=-1.453954865e-08 ppdiblc2=2.757922164e-15 pdiblcb=-1.925435828e+00 lpdiblcb=2.294715811e-07 wpdiblcb=1.024884069e-05 ppdiblcb=-1.287559470e-12 drout=1.866253648e+00 ldrout=-1.658754460e-07 wdrout=-2.632260333e-06 pdrout=5.040410022e-13 pscbe1=8.144649871e+08 lpscbe1=-2.769842528e+00 wpscbe1=-5.155451510e+01 ppscbe1=9.871967878e-6 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.903829784e-06 lalpha0=-7.531177975e-13 walpha0=3.721578344e-11 palpha0=-8.492661530e-19 alpha1=-2.006286042e+00 lalpha1=5.469387891e-07 walpha1=1.589683192e-05 palpha1=-3.044020756e-12 beta0=3.916519703e+01 lbeta0=-3.970185429e-06 wbeta0=-9.039575907e-05 pbeta0=1.824432812e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-5.320928991e-01 lkt1=3.733889775e-08 wkt1=1.291575174e-06 pkt1=-1.862373401e-13 kt2=-1.383569620e-01 lkt2=1.234692268e-08 wkt2=6.446899345e-07 pkt2=-7.784022541e-14 at=3.533271257e+04 lat=-2.407677158e-03 wat=-1.884081679e-01 pat=4.033287382e-8 ute=-8.096008382e-01 lute=-1.204490144e-07 wute=1.122672320e-05 pute=-1.383836330e-12 ua1=3.467186280e-09 lua1=-4.928384357e-16 wua1=1.046881540e-14 pua1=-1.242308253e-21 ub1=-3.608840737e-18 lub1=5.910343365e-25 wub1=-5.733111912e-25 pub1=-2.196285018e-31 uc1=-5.174482148e-11 luc1=3.223755714e-17 wuc1=4.891104978e-16 puc1=-1.293443854e-22 kt1l=0.0 prt=0.0 tvoff=-4.536190362e-03 ltvoff=8.272251382e-10 wtvoff=2.365530433e-08 ptvoff=-3.938842089e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.17 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.841795732e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.785153534e-08 wvth0=2.372881924e-07 pvth0=-3.399787704e-14 k1=8.251290249e-01 lk1=7.342205005e-09 wk1=8.986146222e-08 pk1=-9.925786954e-15 k2=-1.334656553e-01 lk2=5.202784046e-09 wk2=-3.284475759e-07 pk2=3.456938350e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.163202145e+00 ldsub=-9.172051666e-08 wdsub=-3.815287776e-06 pdsub=4.555956453e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=4.832417509e-02 lcdscd=-5.214685748e-09 wcdscd=-1.857426862e-07 pcdscd=2.256513598e-14 cit=0.0 voff='-4.736483521e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.573465875e-08 wvoff=-1.389349413e-06 pvoff=2.219492672e-13 nfactor=2.596904091e+00 lnfactor=5.117445421e-08 wnfactor=7.808422968e-07 pnfactor=-4.251856640e-13 eta0=5.541292930e-02 leta0=-4.982306361e-09 weta0=4.750770502e-07 peta0=-4.357296241e-14 etab=1.549630644e-02 letab=-6.291787900e-09 wetab=-3.211877209e-09 petab=7.159226850e-15 u0=3.923127552e-02 lu0=-1.459584679e-09 wu0=1.555712192e-07 pu0=-1.990602797e-14 ua=4.322858429e-09 lua=-6.184892994e-16 wua=5.924133351e-16 pua=-1.186367247e-23 ub=-4.514066654e-18 lub=7.768324587e-25 wub=1.107896289e-23 pub=-1.691079346e-30 uc=1.515404895e-10 luc=-6.372164490e-18 wuc=2.549860830e-16 puc=-4.180034738e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.321081434e+05 lvsat=-8.699592332e-03 wvsat=-7.952667999e-01 pvsat=7.039852318e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.030511266e-01 lketa=9.424962081e-08 wketa=4.040362787e-06 pketa=-5.010818274e-13 dwg=0.0 dwb=0.0 pclm=-6.423937334e-01 lpclm=8.024712324e-08 wpclm=9.024574248e-06 ppclm=-8.675432921e-13 pdiblc1=5.456656013e-03 lpdiblc1=4.471693312e-08 wpdiblc1=2.340152626e-06 ppdiblc1=-2.831575250e-13 pdiblc2=-3.022559731e-03 lpdiblc2=1.298623078e-09 wpdiblc2=6.774271153e-08 ppdiblc2=-7.238220496e-15 pdiblcb=-4.221910571e-01 lpdiblcb=4.684838684e-08 wpdiblcb=5.091244419e-07 ppdiblcb=-1.043203019e-13 drout=-5.905571939e-02 ldrout=6.802268777e-08 wdrout=9.308251097e-06 pdrout=-9.465639694e-13 pscbe1=8.080977076e+08 lpscbe1=-1.996307203e+00 wpscbe1=2.911495519e+01 ppscbe1=7.175661007e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.748579041e-05 lalpha0=1.602449601e-12 walpha0=1.223976838e-10 palpha0=-1.119767450e-17 alpha1=7.514667432e+00 lalpha1=-6.097237647e-07 walpha1=-3.709260781e-05 palpha1=3.393454318e-12 beta0=-1.600527542e+01 lbeta0=2.732254587e-06 wbeta0=2.420836313e-04 pbeta0=-2.214726309e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-4.447132841e-01 lkt1=2.672349784e-08 wkt1=3.671375924e-07 pkt1=-7.393111611e-14 kt2=-5.703568577e-02 lkt2=2.467526113e-09 wkt2=2.518027652e-09 pkt2=1.746708674e-16 at=1.626598428e+05 lat=-1.787614090e-02 wat=-8.201555523e-01 pat=1.170813366e-7 ute=-7.293472729e+00 lute=6.672506461e-07 wute=-6.648878318e-07 pute=6.082792818e-14 ua1=-9.762492427e-09 lua1=1.114382312e-15 wua1=1.024135287e-14 pua1=-1.214674740e-21 ub1=6.179723408e-18 lub1=-5.981391673e-25 wub1=-5.771021949e-24 pub1=4.118205873e-31 uc1=2.377584475e-10 luc1=-2.933036990e-18 wuc1=-1.326957022e-15 puc1=9.128239330e-23 kt1l=0.0 prt=0.0 tvoff=1.258951866e-02 ltvoff=-1.253308748e-09 wtvoff=-5.908867941e-08 ptvoff=6.113393519e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.18 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.405072541e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.191843650e-08 wvth0=-2.549797516e-09 pvth0=2.548305527e-13 k1=5.438947480e-01 lk1=-3.027325579e-07 wk1=-1.713237114e-08 pk1=1.712234631e-12 k2=-3.227934328e-02 lk2=9.705640341e-08 wk2=5.265710843e-09 pk2=-5.262629665e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.829906714e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.202917375e-06 wvoff=9.937918040e-08 pvoff=-9.932102966e-12 nfactor=1.962474827e+00 lnfactor=7.182946238e-05 wnfactor=2.133891330e-06 pnfactor=-2.132642704e-10 eta0=0.08 etab=-0.07 u0=3.254325208e-02 lu0=5.321676185e-09 wu0=1.349748263e-09 pu0=-1.348958471e-13 ua=-7.606625305e-10 lua=2.655905552e-16 wua=-3.428247179e-17 pua=3.426241174e-21 ub=1.751914081e-18 lub=-1.639967959e-24 wub=6.505858451e-26 pub=-6.502051613e-30 uc=5.896148868e-11 luc=-9.713801421e-16 wuc=-4.572057236e-17 puc=4.569381943e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.305507040e+00 la0=-2.726007940e-06 wa0=-1.398551652e-07 pa0=1.397733303e-11 ags=4.631222040e-01 lags=-7.755663179e-07 wags=-2.654889245e-08 pags=2.653335763e-12 a1=0.0 a2=0.42385546 b0=7.933443285e-25 lb0=-7.928801110e-29 wb0=-3.983089923e-30 pb0=3.980759257e-34 b1=2.632636637e-24 lb1=-5.249868664e-29 keta=-9.245430962e-03 lketa=4.505671623e-08 wketa=-9.999795520e-10 pketa=9.993944240e-14 dwg=0.0 dwb=0.0 pclm=1.621466297e-02 lpclm=1.009542633e-06 wpclm=-1.256753424e-08 ppclm=1.256018047e-12 pdiblc1=0.39 pdiblc2=2.768229290e-03 lpdiblc2=3.050508080e-08 wpdiblc2=1.381978157e-09 ppdiblc2=-1.381169506e-13 pdiblcb=-9.611472864e-01 lpdiblcb=9.355995092e-05 wpdiblcb=4.700051023e-06 ppdiblcb=-4.697300835e-10 drout=0.56 pscbe1=8.069316253e+08 lpscbe1=-5.222688733e+03 wpscbe1=-1.870963165e+02 ppscbe1=1.869868390e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.071614333e-01 lkt1=-5.865132761e-07 wkt1=-1.523452037e-08 pkt1=1.522560604e-12 kt2=-4.358994108e-02 lkt2=-1.722387495e-07 wkt2=-8.407037756e-09 pkt2=8.402118462e-13 at=140000.0 ute=-1.760713718e+00 lute=-5.265545319e-06 wute=-1.765389829e-07 pute=1.764356829e-11 ua1=4.321878083e-10 lua1=-5.613494224e-15 wua1=-1.356741777e-16 pua1=1.355947893e-20 ub1=-6.475928878e-19 lub1=7.968222511e-25 wub1=-1.373942042e-25 pub1=1.373138093e-29 uc1=1.483119541e-11 luc1=9.979333129e-17 wuc1=3.514893041e-18 puc1=-3.512836336e-22 kt1l=0.0 prt=0.0 tvoff=7.428050165e-04 ltvoff=2.262824991e-08 wtvoff=8.014189376e-11 ptvoff=-8.009499953e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.19 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.399095837e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=1.022911739e-8 k1=5.287137050e-01 wk1=6.873056959e-8 k2=-2.741228356e-02 wk2=-2.112464776e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.725216033e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-3.986831489e-7 nfactor=5.564486351e+00 wnfactor=-8.560611098e-6 eta0=0.08 etab=-0.07 u0=3.281011666e-02 wu0=-5.414835234e-9 ua=-7.473440369e-10 wua=1.375322653e-16 ub=1.669675077e-18 wub=-2.609979397e-25 uc=1.024996628e-11 wuc=1.834189182e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.168806699e+00 wa0=5.610621602e-7 ags=4.242301015e-01 wags=1.065071778e-7 a1=0.0 a2=0.42385546 b0=-3.182688907e-24 wb0=1.597910977e-29 b1=0.0 keta=-6.985984688e-03 wketa=4.011655107e-9 dwg=0.0 dwb=0.0 pclm=6.683990892e-02 wpclm=5.041764384e-8 pdiblc1=0.39 pdiblc2=4.297958860e-03 wpdiblc2=-5.544133097e-9 pdiblcb=3.730576837e+00 wpdiblcb=-1.885536925e-5 drout=0.56 pscbe1=5.450309458e+08 wpscbe1=7.505812417e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.365731470e-01 wkt1=6.111689117e-8 kt2=-5.222714843e-02 wkt2=3.372682560e-8 at=140000.0 ute=-2.024763514e+00 wute=7.082279944e-7 ua1=1.506895175e-10 wua1=5.442891375e-16 ub1=-6.076348700e-19 wub1=5.511894316e-25 uc1=1.983550308e-11 wuc1=-1.410082695e-17 kt1l=0.0 prt=0.0 tvoff=1.877537398e-03 wtvoff=-3.215082116e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.20 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.373391674e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.041292537e-08 wvth0=-8.547558013e-09 pvth0=1.491147049e-13 k1=5.140462892e-01 lk1=1.164810769e-07 wk1=1.036439781e-07 pk1=-2.772643450e-13 k2=-1.944187180e-02 lk2=-6.329691336e-08 wk2=-2.690422874e-08 pk2=4.589846149e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.188275770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.264103588e-07 wvoff=-6.344300993e-07 pvoff=1.872181106e-12 nfactor=7.961284143e+00 lnfactor=-1.903413611e-05 wnfactor=-1.585415027e-05 pnfactor=5.792153920e-11 eta0=0.08 etab=-0.07 u0=3.075792336e-02 lu0=1.629746436e-08 wu0=1.690115281e-09 pu0=-5.642386504e-14 ua=-6.370634142e-10 lua=-8.757920210e-16 wua=-3.667156890e-16 pua=4.004478069e-21 ub=1.274733400e-18 lub=3.136423797e-24 wub=1.234560894e-24 pub=-1.187695954e-29 uc=-1.036975530e-10 luc=9.049126293e-16 wuc=5.583472091e-16 puc=-2.977487774e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=8.676959089e-01 la0=2.391267120e-06 wa0=1.978129559e-06 pa0=-1.125362091e-11 ags=2.767219081e-01 lags=1.171434253e-06 wags=4.878851410e-07 pags=-3.028707755e-12 a1=0.0 a2=0.42385546 b0=-6.318819849e-24 lb0=2.490553997e-29 wb0=3.172446914e-29 pb0=-1.250415510e-34 b1=0.0 keta=-9.941787502e-03 lketa=2.347346667e-08 wketa=-1.857525663e-09 pketa=4.661001692e-14 dwg=0.0 dwb=0.0 pclm=-3.525093108e-01 lpclm=3.330255958e-06 wpclm=1.107077329e-07 ppclm=-4.787928983e-13 pdiblc1=0.39 pdiblc2=5.730110479e-03 lpdiblc2=-1.137341204e-08 wpdiblc2=-1.293190981e-08 ppdiblc2=5.866992531e-14 pdiblcb=7.431215218e+00 lpdiblcb=-2.938856789e-05 wpdiblcb=-3.743491272e-05 ppdiblcb=1.475491844e-10 drout=0.56 pscbe1=2.964352856e+08 lpscbe1=1.974218955e+03 wpscbe1=1.482197326e+03 ppscbe1=-5.810118889e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.578352919e-01 lkt1=1.688530260e-07 wkt1=1.319497136e-07 pkt1=-5.625178679e-13 kt2=-6.270065129e-02 lkt2=8.317517632e-08 wkt2=6.863781326e-08 pkt2=-2.772451198e-13 at=140000.0 ute=-2.367789449e+00 lute=2.724135661e-06 wute=1.663126171e-06 pute=-7.583310498e-12 ua1=-4.902935981e-10 lua1=5.090358439e-15 wua1=2.612158871e-15 pua1=-1.642195854e-20 ub1=-1.848345385e-19 lub1=-3.357662913e-24 wub1=-9.474477159e-25 pub1=1.190140593e-29 uc1=2.800686194e-11 luc1=-6.489273201e-17 wuc1=-7.445273784e-17 puc1=4.792838554e-22 kt1l=0.0 prt=0.0 tvoff=3.034587883e-03 ltvoff=-9.188700225e-09 wtvoff=-1.460586670e-09 ptvoff=9.045975629e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.21 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.288978976e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.368407210e-08 wvth0=4.302733159e-08 pvth0=-5.416700046e-14 k1=5.393976669e-01 lk1=1.655897643e-08 wk1=3.394633101e-09 pk1=1.178670449e-13 k2=-2.774209482e-02 lk2=-3.058170054e-08 wk2=-1.757834367e-08 pk2=9.140616049e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.291061505e+00 ldsub=-2.881468689e-06 wdsub=-2.208267777e-06 pdsub=8.703856528e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.277796861e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.022853996e-09 wvoff=-2.501296403e-07 pvoff=3.574662271e-13 nfactor=3.040334834e+00 lnfactor=3.617167006e-07 wnfactor=-2.609037513e-06 pnfactor=5.716112711e-12 eta0=2.737312989e-01 leta0=-7.635892025e-07 weta0=-5.851909610e-07 peta0=2.306521980e-12 etab=-2.393625818e-01 letab=6.675402452e-07 wetab=5.115820343e-07 petab=-2.016393426e-12 u0=3.829612064e-02 lu0=-1.341423471e-08 wu0=-2.234164172e-08 pu0=3.829696873e-14 ua=-8.880921376e-10 lua=1.136341777e-16 wua=1.173842263e-15 pua=-2.067609532e-21 ub=2.439480886e-18 lub=-1.454412114e-24 wub=-3.560610616e-24 pub=7.023141833e-30 uc=1.670334835e-10 luc=-1.621699611e-16 wuc=-3.315147767e-16 puc=5.298907855e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.432191236e+00 la0=-3.775169307e-06 wa0=-4.540418939e-06 pa0=1.443914674e-11 ags=6.128729780e-01 lags=-1.535004832e-07 wags=-1.172512311e-06 pags=3.515725557e-12 a1=0.0 a2=0.42385546 b0=3.089572977e-24 lb0=-1.217750864e-29 wb0=-1.551160896e-29 pb0=6.113878954e-35 b1=0.0 keta=-1.066291862e-02 lketa=2.631579489e-08 wketa=2.698194840e-08 pketa=-6.706036636e-14 dwg=0.0 dwb=0.0 pclm=6.020763159e-01 lpclm=-4.322299260e-07 wpclm=-3.866146677e-07 ppclm=1.481396381e-12 pdiblc1=0.39 pdiblc2=3.453475875e-04 lpdiblc2=9.850555515e-09 wpdiblc2=5.521361156e-09 ppdiblc2=-1.406338384e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.824873369e+08 lpscbe1=5.845159942e+01 wpscbe1=7.735031971e+01 ppscbe1=-2.729340824e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.954561531e-01 lkt1=-7.701347615e-08 wkt1=-5.934938309e-08 pkt1=1.914848436e-13 kt2=-4.018358365e-02 lkt2=-5.575530546e-09 wkt2=-7.580472477e-09 pkt2=2.316818642e-14 at=1.615640480e+05 lat=-8.499439328e-02 wat=7.876155072e-03 pat=-3.104375495e-8 ute=-1.519633573e+00 lute=-6.188588514e-07 wute=-1.255302874e-06 pute=3.919636723e-12 ua1=1.256112563e-09 lua1=-1.793076995e-15 wua1=-3.692073731e-15 pua1=8.426086003e-21 ub1=-1.509057963e-18 lub1=1.861745176e-24 wub1=3.666090790e-24 pub1=-6.282791506e-30 uc1=3.232283294e-12 luc1=3.275592290e-17 wuc1=2.030107823e-17 puc1=1.058130159e-22 kt1l=0.0 prt=0.0 tvoff=1.054736371e-03 ltvoff=-1.385143207e-09 wtvoff=5.895837329e-10 ptvoff=9.652576890e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.22 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.499802494e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.275298115e-08 wvth0=-1.226494517e-08 pvth0=5.318218077e-14 k1=4.339235910e-01 lk1=2.213354181e-07 wk1=5.864866327e-07 pk1=-1.014197909e-12 k2=-7.308673911e-03 lk2=-7.025290117e-08 wk2=-2.004148503e-07 pk2=3.641151340e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.472726068e+00 ldsub=2.484386192e-06 wdsub=6.993282230e-06 pdsub=-9.160823989e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.055355787e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.016376899e-08 wvoff=-4.253784392e-09 pvoff=-1.198983048e-13 nfactor=3.742782505e+00 lnfactor=-1.002075619e-06 wnfactor=1.054679293e-06 pnfactor=-1.396942177e-12 eta0=-2.297118130e-01 leta0=2.138385511e-07 weta0=1.155837454e-06 peta0=-1.073660313e-12 etab=8.385251423e-02 letab=4.002266121e-08 wetab=-4.238510134e-07 petab=-2.002632600e-13 u0=3.576247137e-02 lu0=-8.495190128e-09 wu0=-1.303018276e-09 pu0=-2.549224147e-15 ua=-3.621538779e-10 lua=-9.074675903e-16 wua=6.404160834e-16 pua=-1.031970072e-21 ub=1.252708347e-18 lub=8.496901568e-25 wub=-3.725473979e-25 pub=8.335617283e-31 uc=1.491065762e-10 luc=-1.273651214e-16 wuc=-2.873549317e-16 puc=4.441550646e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.458039179e+04 lvsat=2.993695347e-02 wvsat=5.913270429e-02 pvsat=-1.148053175e-7 a0=-1.057509906e+00 la0=3.000036603e-06 wa0=9.021626616e-06 pa0=-1.189137484e-11 ags=-5.230910516e-01 lags=2.051957777e-06 wags=2.780686106e-06 pags=-4.159353825e-12 a1=0.0 a2=0.42385546 b0=-6.179145955e-24 lb0=5.817579409e-30 wb0=3.102321791e-29 pb0=-2.920792534e-35 b1=0.0 keta=9.074946826e-02 lketa=-1.705749345e-07 wketa=-1.259047076e-07 pketa=2.297669359e-13 dwg=0.0 dwb=0.0 pclm=1.210923210e+00 lpclm=-1.614297647e-06 wpclm=-3.230523508e-06 ppclm=7.002805580e-12 pdiblc1=2.309377685e-01 lpdiblc1=3.088170956e-07 wpdiblc1=-1.752455482e-07 ppdiblc1=3.402367784e-13 pdiblc2=3.250864417e-03 lpdiblc2=4.209535267e-09 wpdiblc2=9.288886174e-09 ppdiblc2=-2.137798092e-14 pdiblcb=-4.858075784e-02 lpdiblcb=4.578171121e-08 wpdiblcb=6.768201901e-10 ppdiblcb=-1.314036924e-15 drout=8.424458000e-01 ldrout=-5.483645665e-7 pscbe1=5.795484661e+08 lpscbe1=4.524545760e+02 wpscbe1=1.698512709e+03 ppscbe1=-3.420398165e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.933706367e-06 lalpha0=1.740291042e-11 walpha0=2.699415447e-11 palpha0=-5.240877298e-17 alpha1=1.083892512e+00 lalpha1=-4.540990378e-07 walpha1=-1.335001292e-06 palpha1=2.591886318e-12 beta0=7.605188726e+00 lbeta0=1.214362852e-05 wbeta0=1.699092553e-05 pbeta0=-3.298764405e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.665670832e-01 lkt1=6.104739905e-08 wkt1=-5.676532187e-08 pkt1=1.864679249e-13 kt2=-7.208669111e-02 lkt2=5.636390595e-08 wkt2=7.559956404e-08 pkt2=-1.383246900e-13 at=1.752160667e+05 lat=-1.114995964e-01 wat=-4.090163561e-02 pat=6.365764276e-8 ute=-3.240900578e+00 lute=2.722956941e-06 wute=3.828089819e-06 pute=-5.949699022e-12 ua1=-2.455125386e-09 lua1=5.412239525e-15 wua1=5.976682819e-15 pua1=-1.034566948e-20 ub1=5.047346025e-19 lub1=-2.048004897e-24 wub1=2.050488121e-25 pub1=4.367730397e-31 uc1=-1.021905984e-10 luc1=2.374329717e-16 wuc1=6.150147580e-16 puc1=-1.048815267e-21 kt1l=0.0 prt=0.0 tvoff=6.429926992e-04 ltvoff=-5.857486333e-10 wtvoff=-4.025890135e-10 ptvoff=2.891547186e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.23 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.379757599e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.405503995e-08 wvth0=1.166017521e-07 pvth0=-6.814401061e-14 k1=9.708711841e-01 lk1=-2.841932235e-07 wk1=-1.590937320e-06 pk1=1.035816258e-12 k2=-1.889288381e-01 lk2=1.007399408e-07 wk2=5.693208542e-07 pk2=-3.605802555e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.845205924e+00 ldsub=-6.394003278e-07 wdsub=-4.974679692e-06 pdsub=2.106844609e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.363352714e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.116628958e-08 wvoff=-2.416455083e-07 pvoff=1.036026798e-13 nfactor=2.180179687e+00 lnfactor=4.690930585e-07 wnfactor=-2.000431052e-06 pnfactor=1.479401441e-12 eta0=-4.375200898e-01 leta0=4.094871344e-07 weta0=2.908893583e-08 peta0=-1.284235793e-14 etab=2.377964480e-01 letab=-1.049133972e-07 wetab=-1.196533814e-06 petab=5.272067793e-13 u0=2.838322382e-02 lu0=-1.547731865e-09 wu0=-3.859644249e-10 pu0=-3.412617509e-15 ua=-1.187563307e-09 lua=-1.303561687e-16 wua=-5.731842773e-16 pua=1.106176777e-22 ub=2.124290389e-18 lub=2.910786637e-26 wub=8.143792299e-25 pub=-2.839130748e-31 uc=-5.360119431e-11 luc=6.348140659e-17 wuc=3.855931819e-16 puc=-1.894161631e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.150570059e+04 lvsat=1.400201219e-02 wvsat=-1.306986695e-01 pvsat=6.391826329e-8 a0=2.684353664e+00 la0=-5.228755617e-07 wa0=-6.795279368e-06 pa0=3.000020707e-12 ags=1.927752772e+00 lags=-2.554773711e-07 wags=-2.643538753e-06 pags=9.474779406e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.690295081e-01 lketa=7.400333490e-08 wketa=3.135728086e-07 pketa=-1.839949929e-13 dwg=0.0 dwb=0.0 pclm=-1.354558376e+00 lpclm=8.010673488e-07 wpclm=8.082443802e-06 ppclm=-3.648194761e-12 pdiblc1=-2.279330893e-01 lpdiblc1=7.408375840e-07 wpdiblc1=2.884591810e-06 ppdiblc1=-2.540557257e-12 pdiblc2=9.345103594e-03 lpdiblc2=-1.528105599e-09 wpdiblc2=-1.248908139e-08 ppdiblc2=-8.743293506e-16 pdiblcb=2.216151568e-02 lpdiblcb=-2.082114891e-08 wpdiblcb=-1.353640380e-09 ppdiblcb=5.976132769e-16 drout=-2.100302390e-01 ldrout=4.425268896e-07 wdrout=-5.538903931e-07 pdrout=5.214800507e-13 pscbe1=1.289805086e+09 lpscbe1=-2.162420883e+02 wpscbe1=-3.642544457e+03 ppscbe1=1.608132382e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.223816197e-05 lalpha0=-1.194496721e-11 walpha0=-7.548037552e-11 palpha0=4.406956236e-17 alpha1=3.822149758e-01 lalpha1=2.065205392e-07 walpha1=2.670002584e-06 palpha1=-1.178768761e-12 beta0=3.191459305e+01 lbeta0=-1.074333532e-05 wbeta0=-6.182110741e-05 pbeta0=4.121278159e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.231224660e-01 lkt1=2.014490020e-08 wkt1=2.705583915e-07 pkt1=-1.217027687e-13 kt2=8.288969881e-03 lkt2=-1.930865361e-08 wkt2=-1.303606866e-07 pkt2=5.558400254e-14 at=4.972053216e+04 lat=6.652692389e-03 wat=9.882949145e-02 pat=-6.789725712e-8 ute=9.345689416e-01 lute=-1.208189155e-06 wute=-6.155521500e-06 pute=3.449731264e-12 ua1=5.301043958e-09 lua1=-1.890085326e-15 wua1=-9.495607175e-15 pua1=4.221274941e-21 ub1=-1.398061313e-18 lub1=-2.565491820e-25 wub1=-2.474547094e-24 pub1=2.959575071e-30 uc1=3.801136189e-10 luc1=-2.166496965e-16 wuc1=-1.373376917e-15 puc1=8.232276573e-22 kt1l=0.0 prt=0.0 tvoff=-1.184977636e-03 ltvoff=1.135259846e-09 wtvoff=4.683567792e-09 ptvoff=-1.896998240e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.24 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.426728896e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.216727702e-08 wvth0=-7.712981251e-08 pvth0=1.738576294e-14 k1=7.509977129e-03 lk1=1.411172624e-07 wk1=1.254092729e-06 pk1=-2.202246776e-13 k2=1.248967557e-01 lk2=-3.780966534e-08 wk2=-4.093691447e-07 pk2=7.149767735e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.301309091e-01 ldsub=2.948408043e-08 wdsub=-5.644007330e-07 pdsub=1.597681924e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.497814002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.230011963e-09 wvoff=-4.409732783e-08 pvoff=1.638792376e-14 nfactor=5.099072746e+00 lnfactor=-8.195573624e-07 wnfactor=-4.579979495e-06 pnfactor=2.618235965e-12 eta0=0.49 etab=1.669882494e-03 letab=-6.668243145e-10 wetab=-6.931995496e-09 petab=2.014230863e-15 u0=2.995991325e-02 lu0=-2.243818172e-09 wu0=-1.154355212e-08 pu0=1.513301253e-15 ua=-9.768703982e-10 lua=-2.233741381e-16 wua=-7.188610272e-16 pua=1.749319232e-22 ub=1.851131692e-18 lub=1.497036068e-25 wub=5.619952383e-25 pub=-1.724890759e-31 uc=1.537169811e-10 luc=-2.804666542e-17 wuc=-2.321205299e-16 puc=8.329579270e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.275121644e+05 lvsat=-6.309197498e-03 wvsat=-6.602797150e-02 pvsat=3.536705550e-8 a0=1.5 ags=2.367433823e+00 lags=-4.495903998e-07 wags=-8.784281852e-07 pags=1.682063365e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.351771810e-02 lketa=-6.588709825e-09 wketa=-1.382023008e-07 pketa=1.545739302e-14 dwg=0.0 dwb=0.0 pclm=3.660302697e-01 lpclm=4.145155021e-08 wpclm=2.846237165e-07 ppclm=-2.055663626e-13 pdiblc1=1.780088717e+00 lpdiblc1=-1.456759311e-07 wpdiblc1=-3.069404975e-06 ppdiblc1=8.804896803e-14 pdiblc2=8.508210237e-03 lpdiblc2=-1.158628898e-09 wpdiblc2=-2.583911049e-08 ppdiblc2=5.019521596e-15 pdiblcb=-2.563634957e-01 lpdiblcb=1.021437442e-07 wpdiblcb=1.161590970e-06 ppdiblcb=-5.128261510e-13 drout=6.332619180e-01 ldrout=7.022520838e-08 wdrout=1.107780786e-06 pdrout=-2.121245116e-13 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.334344912e-05 lalpha0=3.763815942e-12 walpha0=4.995367898e-11 palpha0=-1.130781663e-17 alpha1=0.85 beta0=-1.796772980e+00 lbeta0=4.139760825e-06 wbeta0=5.728731617e-05 pbeta0=-1.137191990e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.489901360e-01 lkt1=-1.258348562e-08 wkt1=-1.672344884e-07 pkt1=7.157665873e-14 kt2=-3.156033119e-02 lkt2=-1.715745077e-09 wkt2=-6.203417111e-08 pkt2=2.541880254e-14 at=8.839446660e+04 lat=-1.042130823e-02 wat=-7.096684773e-02 pat=7.065449474e-9 ute=-2.272617170e+00 lute=2.077386122e-07 wute=8.296971517e-07 pute=3.658550223e-13 ua1=1.321367232e-09 lua1=-1.331137668e-16 wua1=-3.960519759e-15 pua1=1.777611338e-21 ub1=-3.502741847e-18 lub1=6.726378082e-25 wub1=1.083283669e-23 pub1=-2.915448566e-30 uc1=-2.894527208e-10 luc1=7.895446850e-17 wuc1=1.034432690e-15 puc1=-2.397865747e-22 kt1l=0.0 prt=0.0 tvoff=3.449349308e-03 ltvoff=-9.107306193e-10 wtvoff=-5.874313625e-09 ptvoff=2.764158595e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.25 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.541739996e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.436957858e-08 wvth0=9.953280571e-08 pvth0=-1.644265517e-14 k1=5.488890272e-01 lk1=3.745075359e-08 wk1=2.286407609e-08 pk1=1.553837214e-14 k2=-2.127373646e-02 lk2=-9.820062482e-09 wk2=-1.221803117e-07 pk2=1.650503647e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.044564707e-01 ldsub=-6.134262406e-08 wdsub=-9.563002741e-08 pdsub=7.000516509e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-3.375693880e-03 lcdscd=1.680422518e-09 wcdscd=4.405952951e-08 pcdscd=-8.436783069e-15 cit=0.0 voff='-4.623305279e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.547017031e-08 wvoff=8.453094268e-07 pvoff=-1.539210181e-13 nfactor=-1.690114708e+00 lnfactor=4.804769863e-07 wnfactor=2.303027229e-05 pnfactor=-2.668740709e-12 eta0=1.178462252e+00 leta0=-1.318308828e-07 weta0=4.855214603e-07 peta0=-9.297056236e-14 etab=-2.928886499e-02 letab=5.261342407e-09 wetab=3.515103868e-07 petab=-6.662246716e-14 u0=5.597482167e-03 lu0=2.421246305e-09 wu0=-1.030112124e-08 pu0=1.275393133e-15 ua=-5.940123990e-09 lua=7.270194391e-16 wua=6.753007260e-15 pua=-1.255826248e-21 ub=7.237824245e-18 lub=-8.817726034e-25 wub=-1.255818361e-23 pub=2.339841490e-30 uc=-1.779758108e-10 luc=3.546786053e-17 wuc=8.392916990e-16 puc=-1.218646494e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.178439355e+04 lvsat=4.361890433e-03 wvsat=2.389782032e-01 pvsat=-2.303735687e-8 a0=1.5 ags=-2.115963811e+00 lags=4.089174795e-07 wags=-5.185673973e-12 pags=6.299867884e-19 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.656575744e-03 lketa=-4.317467119e-09 wketa=-6.886536973e-08 pketa=2.180341435e-15 dwg=0.0 dwb=0.0 pclm=5.492247522e-01 lpclm=6.372371524e-09 wpclm=-3.423910820e-07 ppclm=-8.550180691e-14 pdiblc1=2.088533172e+00 lpdiblc1=-2.047387260e-07 wpdiblc1=-6.895971963e-06 ppdiblc1=8.207829742e-13 pdiblc2=-1.172868874e-02 lpdiblc2=2.716453940e-09 wpdiblc2=1.269063252e-08 ppdiblc2=-2.358384773e-15 pdiblcb=9.497971606e-01 lpdiblcb=-1.288191352e-07 wpdiblcb=-4.186646065e-06 ppdiblcb=5.112863660e-13 drout=5.565724869e-01 ldrout=8.491016078e-08 wdrout=3.943166814e-06 pdrout=-7.550612405e-13 pscbe1=7.880444351e+08 lpscbe1=2.289323296e+00 wpscbe1=8.109335383e+01 ppscbe1=-1.552824195e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=9.831821059e-06 lalpha0=-6.739238438e-13 walpha0=-2.587743248e-12 palpha0=-1.246869851e-18 alpha1=1.628235406e+00 lalpha1=-1.490211850e-07 walpha1=-2.350762771e-06 palpha1=4.501381600e-13 beta0=1.144785664e+01 lbeta0=1.603599678e-06 wbeta0=4.876280706e-05 pbeta0=-9.739595747e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.300703580e-01 lkt1=2.942241761e-09 wkt1=2.772943392e-07 pkt1=-1.354438835e-14 kt2=-2.997663379e-02 lkt2=-2.019000957e-09 wkt2=1.005521904e-07 pkt2=-5.714209485e-15 at=9.921536163e+04 lat=-1.249335814e-02 wat=-5.091394400e-01 pat=9.096936648e-8 ute=1.282631189e+00 lute=-4.730416752e-07 wute=7.223961297e-07 pute=3.864016658e-13 ua1=4.008276405e-09 lua1=-6.476192567e-16 wua1=7.752201005e-15 pua1=-4.652107098e-22 ub1=-1.524146992e-18 lub1=2.937645940e-25 wub1=-1.103979132e-23 pub1=1.272853480e-30 uc1=2.907230703e-10 luc1=-3.214107305e-17 wuc1=-1.230294759e-15 puc1=1.938770254e-22 kt1l=0.0 prt=0.0 tvoff=-4.744525882e-03 ltvoff=6.582817653e-10 wtvoff=2.470128031e-08 ptvoff=-3.090639585e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.26 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='7.932227400e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.126205386e-08 wvth0=-3.101774205e-07 pvth0=3.333140137e-14 k1=7.462977193e-01 lk1=1.346836122e-08 wk1=4.856444379e-07 pk1=-4.068296290e-14 k2=-2.426932034e-01 lk2=1.707930287e-08 wk2=2.199437473e-07 pk2=-2.505824697e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.196620886e-01 ldsub=-2.446893756e-09 wdsub=4.198164250e-07 pdsub=7.385637371e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.533842624e-02 lcdscd=-1.807941078e-09 wcdscd=-7.033972426e-08 pcdscd=5.461124675e-15 cit=0.0 voff='-1.818182746e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.391858708e-09 wvoff=-7.143081722e-07 pvoff=3.555068558e-14 nfactor=2.894881703e+00 lnfactor=-7.653588768e-08 wnfactor=-7.151936367e-07 pnfactor=2.160009652e-13 eta0=3.755941118e-01 leta0=-3.429364389e-08 weta0=-1.132434840e-06 peta0=1.035884768e-13 etab=1.145639643e-01 letab=-1.221476241e-08 wetab=-5.005941302e-07 petab=3.689630220e-14 u0=1.222856432e-01 lu0=-1.175473163e-08 wu0=-2.614141970e-07 pu0=3.178211626e-14 ua=1.359984090e-08 lua=-1.646812735e-15 wua=-4.598390171e-14 pua=5.150969875e-21 ub=-1.179827650e-17 lub=1.430847132e-24 wub=4.765029993e-23 pub=-4.974646340e-30 uc=4.176827894e-10 luc=-3.689632016e-17 wuc=-1.081216464e-15 puc=1.114502054e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.266143320e+04 lvsat=9.114782394e-03 wvsat=2.060817358e-01 pvsat=-1.904089663e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.994216992e-01 lketa=-5.264036090e-08 wketa=-1.996810761e-06 pketa=2.363987153e-13 dwg=0.0 dwb=0.0 pclm=2.073045450e+00 lpclm=-1.787505098e-07 wpclm=-4.608646609e-06 ppclm=4.327885120e-13 pdiblc1=6.446334942e-01 lpdiblc1=-2.932512979e-08 wpdiblc1=-8.689190615e-07 ppdiblc1=8.858042545e-14 pdiblc2=1.358789011e-02 lpdiblc2=-3.591559583e-10 wpdiblc2=-1.565224447e-08 ppdiblc2=1.084877981e-15 pdiblcb=-6.492614905e-01 lpdiblcb=6.544410411e-08 wpdiblcb=1.649161526e-06 ppdiblcb=-1.976825551e-13 drout=3.745694723e+00 ldrout=-3.025235432e-07 wdrout=-9.794000727e-06 pdrout=9.138122954e-13 pscbe1=8.478439750e+08 lpscbe1=-4.975483608e+00 wpscbe1=-1.704364270e+02 ppscbe1=1.502910500e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.725867298e-05 lalpha0=-1.576182376e-12 walpha0=-5.204148092e-11 palpha0=4.761066923e-18 alpha1=-9.658826141e-01 lalpha1=1.661278368e-07 walpha1=5.485113132e-06 palpha1=-5.018110600e-13 beta0=5.754526766e+01 lbeta0=-3.996590397e-06 wbeta0=-1.271865789e-04 pbeta0=1.163579136e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-5.537720552e-01 lkt1=3.011886615e-08 wkt1=9.146815486e-07 pkt1=-9.097801088e-14 kt2=-9.830225710e-02 lkt2=6.281605715e-09 wkt2=2.097022962e-07 pkt2=-1.897441923e-14 at=-1.851984180e+05 lat=2.205893430e-02 wat=9.263127635e-01 pat=-8.341797991e-8 ute=-1.664919315e+01 lute=1.705423937e-06 wute=4.630674151e-05 pute=-5.151458118e-12 ua1=-1.935024749e-08 lua1=2.190114377e-15 wua1=5.837794275e-14 pua1=-6.615529571e-21 ub1=1.155861664e-17 lub1=-1.295608028e-24 wub1=-3.277646541e-23 pub1=3.913555069e-30 uc1=-2.889274245e-10 luc1=3.827834696e-17 wuc1=1.317338921e-15 puc1=-1.156247997e-22 kt1l=0.0 prt=0.0 tvoff=8.710518346e-04 ltvoff=-2.393230918e-11 wtvoff=-2.545698734e-10 ptvoff=-5.885316972e-17 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.27 nmos lmin=2.0e-05 lmax=0.0001 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.357277245e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.509226603e-07 wvth0=1.188740273e-08 pvth0=-2.370524750e-13 k1=5.343413802e-01 lk1=3.415184830e-07 wk1=1.172483735e-08 pk1=-2.338106798e-13 k2=-2.974941862e-02 lk2=-9.285389777e-08 wk2=-2.376260542e-09 pk2=4.738616634e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.728548903e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.312154291e-07 wvoff=6.876271538e-08 pvoff=-1.371230726e-12 nfactor=-3.052561886e-01 lnfactor=6.053629305e-05 wnfactor=8.983872203e-06 pnfactor=-1.791517618e-10 eta0=0.08 etab=-0.07 u0=3.517337258e-02 lu0=-8.287427487e-08 wu0=-6.594877881e-09 pu0=1.315116649e-13 ua=-8.680732743e-10 lua=3.315475337e-15 wua=2.901658580e-16 pua=-5.786338395e-21 ub=2.070853472e-18 lub=-9.723138982e-24 wub=-8.983399452e-25 pub=1.791423344e-29 uc=5.003267722e-11 luc=4.175612121e-16 wuc=-1.874991873e-17 puc=3.739012419e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.253332997e+00 la0=2.018417439e-06 wa0=1.774341638e-08 pa0=-3.538300894e-13 ags=4.793691463e-01 lags=-3.964197182e-07 wags=-7.562492638e-08 pags=1.508073411e-12 a1=0.0 a2=0.42385546 b0=-5.252836681e-25 lb0=5.249763036e-29 b1=7.952226470e-24 lb1=-1.585792128e-28 wb1=-1.606852328e-29 pb1=3.204302320e-34 keta=-1.615900106e-02 lketa=2.094075598e-07 wketa=1.988337152e-08 pketa=-3.965039749e-13 dwg=0.0 dwb=0.0 pclm=-1.155902651e-01 lpclm=3.970773920e-06 wpclm=3.855666493e-07 ppclm=-7.688771939e-12 pdiblc1=0.39 pdiblc2=2.922243663e-03 lpdiblc2=-9.167228003e-09 wpdiblc2=9.167574132e-10 ppdiblc2=-1.828150512e-14 pdiblcb=5.948353765e-01 lpdiblcb=-6.194726860e-05 wpdiblcb=1.942890293e-22 ppdiblcb=1.332267630e-26 drout=0.56 pscbe1=8.968140358e+08 lpscbe1=-2.059920722e+03 wpscbe1=-4.585980021e+02 ppscbe1=9.145125639e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.835034929e-01 lkt1=-6.548087466e-07 wkt1=-8.669645221e-08 pkt1=1.728856088e-12 kt2=-4.587796177e-02 lkt2=9.604417442e-08 wkt2=-1.495769239e-09 pkt2=2.982786133e-14 at=140000.0 ute=-1.641698966e+00 lute=-2.963325433e-06 wute=-5.360387502e-07 pute=1.068940923e-11 ua1=6.824145494e-10 lua1=-7.010121296e-15 wua1=-8.915170793e-16 pua1=1.777817536e-20 ub1=-1.050949859e-18 lub1=1.247917972e-23 wub1=1.080998771e-24 pub1=-2.155672186e-29 uc1=1.297268203e-11 luc1=4.376458165e-17 wuc1=9.128778041e-18 puc1=-1.820413995e-22 kt1l=0.0 prt=0.0 tvoff=-1.361889670e-03 ltvoff=6.247646965e-08 wtvoff=6.437650015e-09 ptvoff=-1.283763076e-13 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.28 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.543296+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.0344057365 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.30450827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.73044 eta0=0.08 etab=-0.07 u0=0.0310175 ua=-7.0181308e-10 ub=1.58327e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.35455 ags=0.45949 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0017711 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.29 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.345094423e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.977832469e-8 k1=5.483583067e-01 lk1=2.469090016e-8 k2=-2.834869287e-02 lk2=-4.810192719e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.288598150e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.933874537e-07 wvoff=-4.440892099e-22 nfactor=2.712663898e+00 lnfactor=1.411686641e-7 eta0=0.08 etab=-0.07 u0=3.131744708e-02 lu0=-2.382025573e-9 ua=-7.584670440e-10 lua=4.499166616e-16 ub=1.683442867e-18 lub=-7.955214184e-25 uc=8.114694611e-11 luc=-8.080419208e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.522568651e+00 la0=-1.334317761e-6 ags=4.382394782e-01 lags=1.687607211e-7 a1=0.0 a2=0.42385546 b0=4.183773362e-24 lb0=-1.649028413e-29 b1=0.0 keta=-1.055673353e-02 lketa=3.890401793e-8 dwg=0.0 dwb=0.0 pclm=-3.158587910e-01 lpclm=3.171748434e-6 pdiblc1=0.39 pdiblc2=1.448917071e-03 lpdiblc2=8.049650856e-9 pdiblcb=-4.961857729e+00 lpdiblcb=1.945855562e-5 drout=0.56 pscbe1=7.871264144e+08 lpscbe1=5.074105736e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141524753e-01 lkt1=-1.737219702e-8 kt2=-3.997765383e-02 lkt2=-8.608635726e-9 at=140000.0 ute=-1.817200642e+00 lute=2.136310714e-7 ua1=3.744786981e-10 lua1=-3.462384507e-16 ub1=-4.984933079e-19 lub1=5.823754382e-25 uc1=3.358795633e-12 luc1=9.377732624e-17 kt1l=0.0 prt=0.0 tvoff=2.551051103e-03 ltvoff=-6.193970768e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.30 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.431423774e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.575173196e-8 k1=5.405214824e-01 lk1=5.557963332e-8 k2=-3.356152058e-02 lk2=-2.755563975e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.105867411e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.213643889e-7 nfactor=2.176595884e+00 lnfactor=2.254073237e-6 eta0=0.08 etab=-0.07 u0=3.089977388e-02 lu0=-7.357724803e-10 ua=-4.994839710e-10 lua=-5.708614947e-16 ub=1.260717430e-18 lub=8.706449708e-25 uc=5.728334625e-11 luc=1.325385269e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=9.290558192e-01 la0=1.005004755e-6 ags=2.247051008e-01 lags=1.010403480e-6 a1=0.0 a2=0.42385546 b0=-2.045646724e-24 lb0=8.062887923e-30 b1=0.0 keta=-1.730367952e-03 lketa=4.115021555e-09 pketa=-3.469446952e-30 dwg=0.0 dwb=0.0 pclm=4.740849990e-01 lpclm=5.819604485e-8 pdiblc1=0.39 pdiblc2=2.173230347e-03 lpdiblc2=5.194780220e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.080946667e+08 lpscbe1=-3.190501548e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.151041549e-01 lkt1=-1.362116500e-8 kt2=-4.269314869e-02 lkt2=2.094449254e-9 at=1.641715007e+05 lat=-9.527163161e-2 ute=-1.935209808e+00 lute=6.787625481e-7 ua1=3.382738202e-11 lua1=9.964339426e-16 ub1=-2.953746049e-19 lub1=-2.182140860e-25 uc1=9.953088154e-12 luc1=6.778601459e-17 kt1l=0.0 prt=0.0 tvoff=1.249921926e-03 ltvoff=-1.065588329e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.31 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.459198590e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.035929028e-8 k1=6.280838306e-01 lk1=-1.144214397e-7 k2=-7.365732226e-02 lk2=5.028979786e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.069438219e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.985688779e-8 nfactor=4.091940991e+00 lnfactor=-1.464542472e-6 eta0=1.529357436e-01 leta0=-1.416037250e-7 etab=-5.646613875e-02 letab=-2.627580214e-8 u0=3.533109864e-02 lu0=-9.339127472e-9 ua=-1.501399406e-10 lua=-1.249108039e-15 ub=1.129374091e-18 lub=1.125646224e-24 uc=5.397584470e-11 luc=1.967532064e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.415666069e+04 lvsat=-8.070098536e-3 a0=1.929158651e+00 la0=-9.366808915e-7 ags=3.974732892e-01 lags=6.749764612e-7 a1=0.0 a2=0.42385546 b0=4.091293448e-24 lb0=-3.851895503e-30 b1=0.0 keta=4.906789049e-02 lketa=-9.450908604e-08 wketa=-1.127570259e-23 pketa=4.336808690e-29 dwg=0.0 dwb=0.0 pclm=1.414372522e-01 lpclm=7.040269881e-7 pdiblc1=1.729215824e-01 lpdiblc1=4.214547087e-7 pdiblc2=6.326011001e-03 lpdiblc2=-2.867785281e-9 pdiblcb=-4.835669208e-02 lpdiblcb=4.534669069e-8 drout=8.424458000e-01 ldrout=-5.483645665e-7 pscbe1=1.141852219e+09 lpscbe1=-6.798906303e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.885203200e-09 lalpha0=5.264299838e-14 alpha1=6.419315940e-01 lalpha1=4.039618973e-7 beta0=1.323014587e+01 lbeta0=1.222852983e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.853596146e-01 lkt1=1.227788264e-7 kt2=-4.705896047e-02 lkt2=1.057061171e-8 at=1.616753124e+05 lat=-9.042531701e-2 ute=-1.973586381e+00 lute=7.532701261e-7 ua1=-4.765054085e-10 lua1=1.987237911e-15 ub1=5.726173542e-19 lub1=-1.903408323e-24 pub1=7.703719778e-46 uc1=1.014140638e-10 luc1=-1.097841893e-16 puc1=-1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=5.097129705e-04 ltvoff=3.715169938e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.32 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.765775334e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.495519092e-9 k1=4.441809683e-01 lk1=5.872053047e-8 k2=-4.514419294e-04 lk2=-1.863251358e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.983056426e-01 ldsub=5.808437373e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.163335990e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.313205586e-8 nfactor=1.517923890e+00 lnfactor=9.588585914e-7 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=-6.245004514e-23 peta0=-1.734723476e-29 etab=-1.583239050e-01 letab=6.962185877e-8 u0=2.825544777e-02 lu0=-2.677501234e-9 ua=-1.377319714e-09 lua=-9.373546230e-17 ub=2.393895965e-18 lub=-6.488341585e-26 uc=7.405195307e-11 luc=7.739456778e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.823705034e+04 lvsat=3.516257173e-2 a0=4.347319399e-01 la0=4.703009348e-7 ags=1.052591960e+00 lags=5.819140435e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.521917686e-02 lketa=1.309058786e-8 dwg=0.0 dwb=0.0 pclm=1.321187562e+00 lpclm=-4.066914119e-7 pdiblc1=7.270299152e-01 lpdiblc1=-1.002305291e-7 pdiblc2=5.210511433e-03 lpdiblc2=-1.817558055e-9 pdiblcb=2.171338417e-02 lpdiblcb=-2.062330512e-08 wpdiblcb=8.239936511e-24 ppdiblcb=-4.336808690e-30 drout=-3.933992800e-01 ldrout=6.151662745e-7 pscbe1=8.391689559e+07 lpscbe1=3.161406654e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.750110526e-06 lalpha0=2.644549936e-12 walpha0=-6.352747104e-28 palpha0=7.411538288e-34 alpha1=1.266136812e+00 lalpha1=-1.837185766e-7 beta0=1.144831069e+01 lbeta0=2.900425854e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.335523391e-01 lkt1=-2.014559817e-8 kt2=-3.486778889e-02 lkt2=-9.072056564e-10 at=8.243868235e+04 lat=-1.582513911e-2 ute=-1.103256752e+00 lute=-6.613303469e-8 ua1=2.157461034e-09 lua1=-4.926046194e-16 ub1=-2.217276329e-18 lub1=7.232375218e-25 uc1=-7.455180121e-11 luc1=5.588520916e-17 puc1=1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=3.655481450e-04 ltvoff=5.072461586e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.33 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.171385602e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.641160638e-8 k1=4.226855856e-01 lk1=6.821044101e-8 k2=-1.062757987e-02 lk2=-1.413989115e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.432823513e-01 ldsub=8.237638655e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.643801093e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.953174921e-10 nfactor=3.582840548e+00 lnfactor=4.722679570e-8 eta0=0.49 etab=-0.000625 u0=2.613834474e-02 lu0=-1.742829885e-9 ua=-1.214854048e-09 lua=-1.654617797e-16 ub=2.037183895e-18 lub=9.259996889e-26 uc=7.687195999e-11 luc=-4.710478990e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.056531722e+05 lvsat=5.399297777e-3 a0=1.5 ags=2.076624421e+00 lags=-3.939045909e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.223505841e-02 lketa=-1.471438664e-9 dwg=0.0 dwb=0.0 pclm=4.602568145e-01 lpclm=-2.660254000e-8 pdiblc1=7.639421041e-01 lpdiblc1=-1.165267438e-7 pdiblc2=-4.599646146e-05 lpdiblc2=5.031165898e-10 pdiblcb=1.281888000e-01 lpdiblcb=-6.763071056e-08 wpdiblcb=-5.551115123e-23 ppdiblcb=-2.775557562e-29 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.194043360e-06 lalpha0=2.028921317e-14 alpha1=0.85 beta0=1.716856810e+01 lbeta0=3.750122900e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.043542083e-01 lkt1=1.111243587e-8 kt2=-5.209714968e-02 lkt2=6.699315923e-9 at=6.490042703e+04 lat=-8.082244924e-3 ute=-1.997940496e+00 lute=3.288573126e-7 ua1=1.021123587e-11 lua1=4.553761050e-16 ub1=8.353966276e-20 lub1=-2.925405273e-25 uc1=5.300299360e-11 luc1=-4.284469763e-19 kt1l=0.0 prt=0.0 tvoff=1.504619322e-03 ltvoff=4.362180831e-12 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.34 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.222536860e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.090611864e-08 wvth0=8.000787264e-07 pvth0=-1.532038750e-13 k1=5.564583292e-01 lk1=4.259483342e-8 k2=3.598162093e-02 lk2=-2.306490057e-08 wk2=-2.951276764e-07 pk2=5.651281824e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=7.727802003e-01 ldsub=-3.816363857e-08 wdsub=5.232872910e-11 pdsub=-1.002021902e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.121050183e-02 lcdscd=-1.112629753e-9 cit=0.0 voff='-1.260427872e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.629434296e-08 wvoff=-1.704920840e-07 pvoff=3.264684719e-14 nfactor=6.043410580e+00 lnfactor=-4.239379174e-07 wnfactor=-3.298616648e-07 pnfactor=6.316389074e-14 eta0=1.339197306e+00 leta0=-1.626093953e-07 weta0=1.292329088e-14 peta0=-2.474628946e-21 etab=1.122004141e-01 letab=-2.160448724e-08 wetab=-7.587665719e-08 petab=1.452931758e-14 u0=-1.334335874e-03 lu0=3.517803835e-09 wu0=1.063735015e-08 pu0=-2.036903631e-15 ua=-3.316293518e-09 lua=2.369344588e-16 wua=-1.172619025e-15 pua=2.245401266e-22 ub=2.430440495e-18 lub=1.729683556e-26 wub=1.963153584e-24 pub=-3.759164272e-31 uc=1.794858784e-10 luc=-2.012017668e-17 wuc=-2.404685181e-16 puc=4.604635465e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.767836467e+05 lvsat=-8.221192264e-03 wvsat=-7.818590070e-02 pvsat=1.497150538e-8 a0=1.5 ags=-2.115965528e+00 lags=4.089176881e-07 wags=-7.216449660e-22 pags=6.245004514e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.213804809e-01 lketa=-5.003526382e-08 wketa=-7.325704288e-07 pketa=1.402769811e-13 dwg=0.0 dwb=0.0 pclm=7.772081259e-02 lpclm=4.664774886e-08 wpclm=1.081848806e-06 ppclm=-2.071589005e-13 pdiblc1=-1.944234950e-01 lpdiblc1=6.698685133e-8 pdiblc2=-7.527371761e-03 lpdiblc2=1.935695220e-09 ppdiblc2=-8.673617380e-31 pdiblcb=-4.362194298e-01 lpdiblcb=4.044556373e-8 drout=1.861983677e+00 ldrout=-1.650578064e-7 pscbe1=8.148909208e+08 lpscbe1=-2.851402867e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=8.975131714e-06 lalpha0=-1.086708271e-12 alpha1=0.85 beta0=2.622343725e+01 lbeta0=-1.358868383e-06 wbeta0=4.131215455e-06 pbeta0=-7.910699226e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.032018945e-01 lkt1=-8.256816093e-09 wkt1=-1.059286014e-07 pkt1=2.028384417e-14 kt2=3.311827170e-03 lkt2=-3.910727419e-9 at=-1.219411189e+05 lat=2.769529534e-02 wat=1.588929021e-01 pat=-3.042576625e-8 ute=1.521785158e+00 lute=-3.451208739e-07 pute=-2.220446049e-28 ua1=6.574693302e-09 lua1=-8.016303080e-16 ub1=-5.178942186e-18 lub1=7.151510720e-25 uc1=-1.165740644e-10 luc1=3.204318556e-17 puc1=1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=3.921987856e-03 ltvoff=-4.585300502e-10 wtvoff=-1.477068418e-09 ptvoff=2.828379231e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.35 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.345917298e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.130607891e-08 wvth0=-1.979664288e-06 pvth0=1.844959848e-13 k1=0.90707349 k2=-3.722707077e-01 lk2=2.653204183e-08 wk2=6.113497036e-07 pk2=-5.361149274e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586854868e-01 ldsub=-5.528208133e-12 wdsub=-1.221003679e-10 pdsub=1.117047426e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-6.697212480e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.975497853e-08 wvoff=7.594671621e-07 pvoff=-8.033018177e-14 nfactor=2.678807818e+00 lnfactor=-1.518578631e-08 wnfactor=-6.251394586e-08 pnfactor=3.068488576e-14 eta0=6.941537032e-04 leta0=-1.365265976e-15 weta0=-3.015434187e-14 peta0=2.758700120e-21 etab=-6.563478702e-02 wetab=4.371998422e-8 u0=5.828081392e-02 lu0=-3.724602253e-09 wu0=-6.807916147e-08 pu0=7.526050500e-15 ua=-2.819282921e-09 lua=1.765546293e-16 wua=3.612229109e-15 pua=-3.567519338e-22 ub=7.944495969e-18 lub=-6.525837078e-25 wub=-1.198535036e-23 pub=1.318631523e-30 uc=1.386863297e-11 wuc=1.385574985e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.921471684e+04 lvsat=8.491506744e-03 wvsat=1.862866775e-01 pvsat=-1.715821025e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.275207956e-01 lketa=7.739155665e-08 wketa=1.709331000e-06 pketa=-1.563798559e-13 dwg=0.0 dwb=0.0 pclm=1.343699992e+00 lpclm=-1.071509977e-07 wpclm=-2.405562380e-06 ppclm=2.165127348e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.863053849e+01 lbeta0=-4.364374842e-07 wbeta0=-9.639502728e-06 pbeta0=8.818795466e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.711670600e-01 wkt1=6.103585679e-8 kt2=-0.028878939 at=2.442027366e+05 lat=-1.678605708e-02 wat=-3.707501049e-01 pat=3.391844410e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=1.227140865e-03 ltvoff=-1.311438687e-10 wtvoff=-1.330183794e-09 ptvoff=2.649934976e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.36 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.416107367e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.360665466e-8 k1=5.401439397e-01 lk1=2.258068246e-7 k2=-3.092541729e-02 lk2=-6.940273678e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.388245892e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.309830202e-6 nfactor=4.140814250e+00 lnfactor=-2.812495837e-5 eta0=0.08 etab=-0.07 u0=3.190960269e-02 lu0=-1.778985329e-8 ua=-7.244717387e-10 lua=4.518473262e-16 ub=1.626269824e-18 lub=-8.574803953e-25 wub=-3.081487911e-39 uc=4.075344244e-11 luc=6.026029425e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.262114120e+00 la0=1.843308815e-6 ags=4.419427736e-01 lags=3.499177697e-7 a1=0.0 a2=0.42385546 b0=-5.252836681e-25 lb0=5.249763036e-29 b1=0.0 keta=-6.318826539e-03 lketa=1.317985732e-8 dwg=0.0 dwb=0.0 pclm=7.522461324e-02 lpclm=1.656416952e-7 pdiblc1=0.39 pdiblc2=3.375942017e-03 lpdiblc2=-1.821464739e-8 pdiblcb=5.948353765e-01 lpdiblcb=-6.194726860e-05 wpdiblcb=2.220446049e-22 ppdiblcb=-2.486899575e-26 drout=0.56 pscbe1=6.698563305e+08 lpscbe1=2.465953182e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.264091047e-01 lkt1=2.007929107e-7 kt2=-4.661820999e-02 lkt2=1.108058239e-7 at=140000.0 ute=-1.906981685e+00 lute=2.326806186e-6 ua1=2.412075017e-10 lua1=1.788202870e-15 ub1=-5.159693327e-19 lub1=1.810873037e-24 uc1=1.749046560e-11 luc1=-4.632673608e-17 kt1l=0.0 prt=0.0 tvoff=1.824068988e-03 ltvoff=-1.056280324e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.37 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.543296+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.0344057365 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.30450827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.73044 eta0=0.08 etab=-0.07 u0=0.0310175 ua=-7.0181308e-10 ub=1.58327e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.35455 ags=0.45949 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0017711 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.38 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.345094423e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.977832469e-8 k1=5.483583067e-01 lk1=2.469090016e-8 k2=-2.834869287e-02 lk2=-4.810192719e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.288598150e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.933874537e-7 nfactor=2.712663898e+00 lnfactor=1.411686641e-7 eta0=0.08 etab=-0.07 u0=3.131744708e-02 lu0=-2.382025573e-9 ua=-7.584670440e-10 lua=4.499166616e-16 ub=1.683442867e-18 lub=-7.955214184e-25 uc=8.114694611e-11 luc=-8.080419208e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.522568651e+00 la0=-1.334317761e-6 ags=4.382394782e-01 lags=1.687607211e-7 a1=0.0 a2=0.42385546 b0=4.183773362e-24 lb0=-1.649028413e-29 b1=0.0 keta=-1.055673353e-02 lketa=3.890401793e-8 dwg=0.0 dwb=0.0 pclm=-3.158587910e-01 lpclm=3.171748434e-06 wpclm=2.220446049e-22 ppclm=-3.552713679e-27 pdiblc1=0.39 pdiblc2=1.448917071e-03 lpdiblc2=8.049650856e-9 pdiblcb=-4.961857729e+00 lpdiblcb=1.945855562e-5 drout=0.56 pscbe1=7.871264144e+08 lpscbe1=5.074105736e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141524753e-01 lkt1=-1.737219702e-8 kt2=-3.997765383e-02 lkt2=-8.608635726e-9 at=140000.0 ute=-1.817200642e+00 lute=2.136310714e-7 ua1=3.744786981e-10 lua1=-3.462384507e-16 ub1=-4.984933079e-19 lub1=5.823754382e-25 uc1=3.358795633e-12 luc1=9.377732624e-17 kt1l=0.0 prt=0.0 tvoff=2.551051103e-03 ltvoff=-6.193970768e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.39 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.431423774e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.575173196e-8 k1=5.405214824e-01 lk1=5.557963332e-8 k2=-3.356152058e-02 lk2=-2.755563975e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.105867411e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.213643889e-7 nfactor=2.176595884e+00 lnfactor=2.254073237e-6 eta0=0.08 etab=-0.07 u0=3.089977388e-02 lu0=-7.357724803e-10 ua=-4.994839710e-10 lua=-5.708614947e-16 ub=1.260717430e-18 lub=8.706449708e-25 uc=5.728334625e-11 luc=1.325385269e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=9.290558192e-01 la0=1.005004755e-6 ags=2.247051008e-01 lags=1.010403480e-6 a1=0.0 a2=0.42385546 b0=-2.045646724e-24 lb0=8.062887923e-30 b1=0.0 keta=-1.730367952e-03 lketa=4.115021555e-09 wketa=1.734723476e-24 pketa=3.469446952e-30 dwg=0.0 dwb=0.0 pclm=4.740849990e-01 lpclm=5.819604485e-8 pdiblc1=0.39 pdiblc2=2.173230347e-03 lpdiblc2=5.194780220e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.080946667e+08 lpscbe1=-3.190501548e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.151041549e-01 lkt1=-1.362116500e-8 kt2=-4.269314869e-02 lkt2=2.094449254e-9 at=1.641715007e+05 lat=-9.527163161e-2 ute=-1.935209808e+00 lute=6.787625481e-7 ua1=3.382738202e-11 lua1=9.964339426e-16 ub1=-2.953746049e-19 lub1=-2.182140860e-25 uc1=9.953088154e-12 luc1=6.778601459e-17 kt1l=0.0 prt=0.0 tvoff=1.249921926e-03 ltvoff=-1.065588329e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.40 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.459198590e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.035929028e-8 k1=6.280838306e-01 lk1=-1.144214397e-7 k2=-7.365732226e-02 lk2=5.028979786e-08 pk2=1.110223025e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.069438219e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.985688779e-8 nfactor=4.091940991e+00 lnfactor=-1.464542472e-6 eta0=1.529357436e-01 leta0=-1.416037250e-7 etab=-5.646613875e-02 letab=-2.627580214e-8 u0=3.533109864e-02 lu0=-9.339127472e-9 ua=-1.501399406e-10 lua=-1.249108039e-15 ub=1.129374091e-18 lub=1.125646224e-24 uc=5.397584470e-11 luc=1.967532064e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.415666069e+04 lvsat=-8.070098536e-3 a0=1.929158651e+00 la0=-9.366808915e-07 wa0=3.552713679e-21 ags=3.974732892e-01 lags=6.749764612e-7 a1=0.0 a2=0.42385546 b0=4.091293448e-24 lb0=-3.851895503e-30 b1=0.0 keta=4.906789049e-02 lketa=-9.450908604e-08 wketa=-1.387778781e-23 pketa=-7.025630078e-29 dwg=0.0 dwb=0.0 pclm=1.414372522e-01 lpclm=7.040269881e-7 pdiblc1=1.729215824e-01 lpdiblc1=4.214547087e-7 pdiblc2=6.326011001e-03 lpdiblc2=-2.867785281e-09 wpdiblc2=1.387778781e-23 pdiblcb=-4.835669208e-02 lpdiblcb=4.534669069e-8 drout=8.424458000e-01 ldrout=-5.483645665e-7 pscbe1=1.141852219e+09 lpscbe1=-6.798906303e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.885203200e-09 lalpha0=5.264299838e-14 alpha1=6.419315940e-01 lalpha1=4.039618973e-7 beta0=1.323014587e+01 lbeta0=1.222852983e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.853596146e-01 lkt1=1.227788264e-7 kt2=-4.705896047e-02 lkt2=1.057061171e-08 wkt2=1.110223025e-22 at=1.616753124e+05 lat=-9.042531701e-2 ute=-1.973586381e+00 lute=7.532701261e-7 ua1=-4.765054085e-10 lua1=1.987237911e-15 ub1=5.726173542e-19 lub1=-1.903408323e-24 uc1=1.014140638e-10 luc1=-1.097841893e-16 puc1=1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=5.097129705e-04 ltvoff=3.715169938e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.41 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.765775334e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.495519092e-9 k1=4.441809683e-01 lk1=5.872053047e-8 k2=-4.514419294e-04 lk2=-1.863251358e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.983056426e-01 ldsub=5.808437373e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.163335990e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.313205586e-8 nfactor=1.517923890e+00 lnfactor=9.588585914e-7 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=2.775557562e-23 peta0=3.955169525e-28 etab=-1.583239050e-01 letab=6.962185877e-8 u0=2.825544777e-02 lu0=-2.677501234e-9 ua=-1.377319714e-09 lua=-9.373546230e-17 ub=2.393895965e-18 lub=-6.488341585e-26 uc=7.405195307e-11 luc=7.739456778e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.823705034e+04 lvsat=3.516257173e-2 a0=4.347319399e-01 la0=4.703009348e-7 ags=1.052591960e+00 lags=5.819140435e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.521917686e-02 lketa=1.309058786e-8 dwg=0.0 dwb=0.0 pclm=1.321187562e+00 lpclm=-4.066914119e-7 pdiblc1=7.270299152e-01 lpdiblc1=-1.002305291e-7 pdiblc2=5.210511433e-03 lpdiblc2=-1.817558055e-9 pdiblcb=2.171338417e-02 lpdiblcb=-2.062330512e-08 wpdiblcb=1.301042607e-23 ppdiblcb=4.553649124e-30 drout=-3.933992800e-01 ldrout=6.151662745e-7 pscbe1=8.391689559e+07 lpscbe1=3.161406654e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.750110526e-06 lalpha0=2.644549936e-12 walpha0=8.470329473e-28 palpha0=1.058791184e-33 alpha1=1.266136812e+00 lalpha1=-1.837185766e-7 beta0=1.144831069e+01 lbeta0=2.900425854e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.335523391e-01 lkt1=-2.014559817e-8 kt2=-3.486778889e-02 lkt2=-9.072056564e-10 at=8.243868235e+04 lat=-1.582513911e-2 ute=-1.103256752e+00 lute=-6.613303469e-8 ua1=2.157461034e-09 lua1=-4.926046194e-16 ub1=-2.217276329e-18 lub1=7.232375218e-25 pub1=1.540743956e-45 uc1=-7.455180121e-11 luc1=5.588520916e-17 wuc1=-5.169878828e-32 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=3.655481450e-04 ltvoff=5.072461586e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.42 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.171385602e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.641160638e-8 k1=4.226855856e-01 lk1=6.821044101e-8 k2=-1.062757987e-02 lk2=-1.413989115e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.432823513e-01 ldsub=8.237638655e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.643801093e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.953174921e-10 nfactor=3.582840548e+00 lnfactor=4.722679570e-8 eta0=0.49 etab=-0.000625 u0=2.613834474e-02 lu0=-1.742829885e-9 ua=-1.214854048e-09 lua=-1.654617797e-16 ub=2.037183895e-18 lub=9.259996889e-26 uc=7.687195999e-11 luc=-4.710478990e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.056531722e+05 lvsat=5.399297777e-3 a0=1.5 ags=2.076624421e+00 lags=-3.939045909e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.223505841e-02 lketa=-1.471438664e-9 dwg=0.0 dwb=0.0 pclm=4.602568145e-01 lpclm=-2.660254000e-8 pdiblc1=7.639421041e-01 lpdiblc1=-1.165267438e-07 ppdiblc1=-2.220446049e-28 pdiblc2=-4.599646146e-05 lpdiblc2=5.031165898e-10 pdiblcb=1.281888000e-01 lpdiblcb=-6.763071056e-8 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.194043360e-06 lalpha0=2.028921317e-14 alpha1=0.85 beta0=1.716856810e+01 lbeta0=3.750122900e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.043542083e-01 lkt1=1.111243587e-8 kt2=-5.209714968e-02 lkt2=6.699315923e-9 at=6.490042703e+04 lat=-8.082244924e-3 ute=-1.997940496e+00 lute=3.288573126e-7 ua1=1.021123587e-11 lua1=4.553761050e-16 ub1=8.353966276e-20 lub1=-2.925405273e-25 uc1=5.300299360e-11 luc1=-4.284469763e-19 kt1l=0.0 prt=0.0 tvoff=1.504619322e-03 ltvoff=4.362180831e-12 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.43 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='7.363788435e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.924445127e-08 wvth0=1.653473812e-07 pvth0=-3.166170864e-14 k1=5.564583292e-01 lk1=4.259483342e-8 k2=-1.444416841e-01 lk2=1.148363641e-08 wk2=6.944142723e-08 pk2=-1.329706113e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=7.728060975e-01 ldsub=-3.816859752e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.121050183e-02 lcdscd=-1.112629753e-9 cit=0.0 voff='-6.763177097e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.747923481e-08 wvoff=-2.885192525e-07 pvoff=5.524739759e-14 nfactor=5.195606966e+00 lnfactor=-2.615953946e-07 wnfactor=1.383237447e-06 pnfactor=-2.648706059e-13 eta0=1.339197312e+00 leta0=-1.626093965e-7 etab=7.464946111e-02 letab=-1.441400546e-08 wetab=-4.857225733e-23 petab=-6.071532166e-30 u0=8.116509315e-03 lu0=1.708099293e-09 wu0=-8.459330064e-09 pu0=1.619843277e-15 ua=-2.676920975e-09 lua=1.145035680e-16 wua=-2.464555646e-15 pua=4.719279024e-22 ub=2.019046042e-18 lub=9.607311382e-26 wub=2.794430381e-24 pub=-5.350942959e-31 uc=-1.068045584e-10 luc=3.470043390e-17 wuc=3.380190998e-16 puc=-6.472592533e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.977280249e+05 lvsat=-1.223174748e-02 wvsat=-1.205067817e-01 pvsat=2.307536159e-8 a0=1.5 ags=-2.115965528e+00 lags=4.089176881e-07 wags=-7.771561172e-22 pags=6.938893904e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.110403275e-01 lketa=5.191586709e-08 wketa=3.432560941e-07 pketa=-6.572873644e-14 dwg=0.0 dwb=0.0 pclm=5.000437792e-01 lpclm=-3.422118672e-08 wpclm=2.284895056e-07 ppclm=-4.375254147e-14 pdiblc1=-1.944234950e-01 lpdiblc1=6.698685133e-8 pdiblc2=-7.527371761e-03 lpdiblc2=1.935695220e-09 ppdiblc2=1.734723476e-30 pdiblcb=-4.362194298e-01 lpdiblcb=4.044556373e-8 drout=1.861983677e+00 ldrout=-1.650578064e-7 pscbe1=8.148909208e+08 lpscbe1=-2.851402867e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=8.975131714e-06 lalpha0=-1.086708271e-12 alpha1=0.85 beta0=2.789901985e+01 lbeta0=-1.679718993e-06 wbeta0=7.454796267e-07 pbeta0=-1.427489118e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-7.115844873e-02 lkt1=-3.354128735e-08 wkt1=-3.727398134e-07 pkt1=7.137445590e-14 kt2=3.311827170e-03 lkt2=-3.910727419e-9 at=-4.330586910e+04 lat=1.263774590e-2 ute=1.521785158e+00 lute=-3.451208739e-07 wute=-1.776356839e-21 pute=2.220446049e-28 ua1=6.574693302e-09 lua1=-8.016303080e-16 ub1=-5.178942186e-18 lub1=7.151510720e-25 wub1=-6.162975822e-39 pub1=7.703719778e-46 uc1=-1.165740644e-10 luc1=3.204318556e-17 kt1l=0.0 prt=0.0 tvoff=4.199106432e-03 ltvoff=-5.115943778e-10 wtvoff=-2.037023080e-09 ptvoff=3.900614015e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.44 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.133420222e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=-9.527284366e-8 k1=0.90707349 k2=-4.991526615e-02 wk2=-4.001201707e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-3.761383875e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=1.662442395e-7 nfactor=3.042310335e+00 wnfactor=-7.970187620e-7 eta0=0.00069413878 etab=-0.043998 u0=2.217655980e-02 wu0=4.874249745e-9 ua=-1.734396174e-09 wua=1.420072232e-15 ub=2.809862381e-18 wub=-1.610145421e-24 uc=1.788286331e-10 wuc=-1.947659564e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.704360465e+04 wvsat=6.943577627e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.163000006e-01 wketa=-1.977835025e-7 dwg=0.0 dwb=0.0 pclm=2.183554635e-01 wpclm=-1.316552145e-7 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.407257900e+01 wbeta0=-4.295439299e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.472502400e-01 wkt1=2.147719650e-7 kt2=-0.028878939 at=60720.487 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-1.203211750e-05 wtvoff=1.173728789e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.45 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.349305493e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.901483927e-07 wvth0=1.136054047e-08 pvth0=-4.362830891e-13 k1=4.463702342e-01 lk1=6.835557268e-06 wk1=1.594745644e-07 pk1=-1.124075312e-11 k2=2.623989744e-03 lk2=-2.573426397e-06 wk2=-5.705519519e-08 pk2=4.258422766e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-5.434008446e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.725271732e-06 wvoff=-3.137402522e-07 pvoff=4.107777159e-12 nfactor=8.411570378e+00 lnfactor=-1.109182155e-04 wnfactor=-7.262984535e-06 pnfactor=1.408008625e-10 eta0=0.08 etab=-0.07 u0=3.344831136e-02 lu0=4.603983980e-08 wu0=-2.616777202e-09 pu0=-1.085508186e-13 ua=-7.622390806e-10 lua=-1.300752883e-15 wua=6.422835002e-17 pua=2.980527999e-21 ub=1.700012982e-18 lub=2.261461885e-24 wub=-1.254099740e-25 pub=-5.304173049e-30 uc=-8.572045330e-11 luc=5.871382155e-15 wuc=2.150855543e-16 puc=-8.960254530e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=9.676267919e-01 la0=8.726934446e-06 wa0=5.008145730e-07 pa0=-1.170651402e-11 ags=3.035505599e-01 lags=9.900747987e-06 wags=2.353542271e-07 pags=-1.624244749e-11 a1=0.0 a2=0.42385546 b0=-1.015401215e-23 lb0=3.726411797e-28 wb0=1.637492378e-29 pb0=-5.444463646e-34 b1=0.0 keta=-5.199211929e-03 lketa=-2.599358382e-07 wketa=-1.904052433e-09 pketa=4.644692916e-13 dwg=0.0 dwb=0.0 pclm=4.989741162e-02 lpclm=6.707037318e-07 wpclm=4.307224956e-08 ppclm=-8.589246615e-13 pdiblc1=0.39 pdiblc2=6.683815899e-03 lpdiblc2=-1.260017528e-07 wpdiblc2=-5.625476174e-09 ppdiblc2=1.833062007e-13 pdiblcb=1.028953664e+01 lpdiblcb=-2.730935842e-04 wpdiblcb=-1.648711919e-05 ppdiblcb=3.590821809e-10 drout=0.56 pscbe1=2.684802298e+08 lpscbe1=1.241583938e+04 wpscbe1=6.825930409e+02 ppscbe1=-1.692109486e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.389762408e-01 lkt1=-9.993845865e-07 wkt1=2.137207380e-08 pkt1=2.041060257e-12 kt2=-4.803677017e-02 lkt2=-1.102829385e-06 wkt2=2.412448837e-09 pkt2=2.063946873e-12 at=140000.0 ute=-1.880757083e+00 lute=-2.875627178e-05 wute=-4.459839711e-08 pute=5.286087705e-11 ua1=7.451040520e-10 lua1=-7.044577113e-14 wua1=-8.569425981e-16 pua1=1.228434077e-19 ub1=-1.185728462e-18 lub1=4.659648383e-23 wub1=1.139013808e-24 pub1=-7.616384286e-29 uc1=-5.505518591e-12 luc1=2.818607852e-15 wuc1=3.910770658e-17 puc1=-4.872199439e-21 kt1l=0.0 prt=0.0 tvoff=2.544595313e-03 ltvoff=-6.014603191e-08 wtvoff=-1.225350126e-09 ptvoff=1.004899224e-13 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.46 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.494805378e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=-1.051762293e-8 k1=7.891509712e-01 wk1=-4.042122700e-7 k2=-1.264248884e-01 wk2=1.564907144e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.411502214e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.077487248e-7 nfactor=2.849386320e+00 wnfactor=-2.022839178e-7 eta0=0.08 etab=-0.07 u0=3.575705805e-02 wu0=-8.060244085e-9 ua=-8.274675637e-10 wua=2.136920359e-16 ub=1.813417865e-18 wub=-3.913968242e-25 uc=2.087100698e-10 wuc=-2.342417692e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.405253880e+00 wa0=-8.622864056e-8 ags=8.000405400e-01 wags=-5.791511460e-7 a1=0.0 a2=0.42385546 b0=8.532718604e-24 wb0=-1.092727249e-29 b1=0.0 keta=-1.823414013e-02 wketa=2.138755641e-8 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=3.652420048e-04 wpdiblc2=3.566727492e-9 pdiblcb=-3.405209289e+00 wpdiblcb=1.519672322e-6 drout=0.56 pscbe1=8.910937792e+08 wpscbe1=-1.659442679e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.890920941e-01 wkt1=1.237245393e-7 kt2=-1.033400402e-01 wkt2=1.059126029e-7 at=140000.0 ute=-3.322789627e+00 wute=2.606200899e-6 ua1=-2.787519902e-09 wua1=5.303250663e-15 ub1=1.150932097e-18 wub1=-2.680352655e-24 uc1=1.358384039e-10 wuc1=-2.052170864e-16 kt1l=0.0 prt=0.0 tvoff=-4.715305619e-04 wtvoff=3.813889298e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.47 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.322720110e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.366612750e-07 wvth0=3.805047358e-09 pvth0=-1.137432855e-13 k1=8.268491944e-01 lk1=-2.993799119e-07 wk1=-4.736105153e-07 pk1=5.511251933e-13 k2=-1.316923254e-01 lk2=4.183127717e-08 wk2=1.757494885e-07 pk2=-1.529432852e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.232062413e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.516467332e-07 wvoff=-9.614648269e-09 pvoff=-7.793303951e-13 nfactor=2.921805899e+00 lnfactor=-5.751190774e-07 wnfactor=-3.556735799e-07 pnfactor=1.218141854e-12 eta0=0.08 etab=-0.07 u0=3.454152540e-02 lu0=9.653135547e-09 wu0=-5.482970748e-09 pu0=-2.046738013e-14 ua=-1.167194515e-09 lua=2.697936825e-15 wua=6.950950158e-16 pua=-3.823055026e-21 ub=2.217347674e-18 lub=-3.207802920e-24 wub=-9.079755997e-25 pub=4.102403114e-30 uc=2.486417791e-10 luc=-3.171171099e-16 wuc=-2.848470728e-16 puc=4.018813100e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.676634318e+00 la0=-2.155163948e-06 wa0=-2.620090035e-07 pa0=1.395957291e-12 ags=7.227959864e-01 lags=6.134365413e-07 wags=-4.839259036e-07 pags=-7.562299295e-13 a1=0.0 a2=0.42385546 b0=1.694061633e-23 lb0=-6.677120211e-29 wb0=-2.169469538e-29 pb0=8.550933810e-35 b1=0.0 keta=-4.138790998e-03 lketa=-1.119380178e-07 wketa=-1.091455845e-08 pketa=2.565267929e-13 dwg=0.0 dwb=0.0 pclm=-1.827285230e-01 lpclm=2.114496274e-06 wpclm=-2.264055939e-07 ppclm=1.797996854e-12 pdiblc1=0.39 pdiblc2=-3.155346759e-03 lpdiblc2=2.795870638e-08 wpdiblc2=7.830158406e-09 ppdiblc2=-3.385797691e-14 pdiblcb=-6.735971186e+00 lpdiblcb=2.645119898e-05 wpdiblcb=3.017114117e-06 ppdiblcb=-1.189191305e-11 drout=0.56 pscbe1=8.162929421e+08 lpscbe1=5.940298001e+02 wpscbe1=-4.960153038e+01 ppscbe1=-9.239342211e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.839300949e-01 lkt1=-4.099394466e-08 wkt1=1.186660528e-07 pkt1=4.017189993e-14 kt2=-9.913620788e-02 lkt2=-3.338467557e-08 wkt2=1.006069301e-07 pkt2=4.213492619e-14 at=140000.0 ute=-2.824199773e+00 lute=-3.959544345e-06 wute=1.712534946e-06 pute=7.097035654e-12 ua1=-2.304822818e-09 lua1=-3.833332137e-15 wua1=4.556505896e-15 pua1=5.930263109e-21 ub1=8.353383867e-19 lub1=2.506283033e-24 wub1=-2.268356862e-24 pub1=-3.271858822e-30 uc1=1.064223906e-10 luc1=2.336068579e-16 wuc1=-1.752732477e-16 puc1=-2.377985761e-22 kt1l=0.0 prt=0.0 tvoff=8.757639968e-04 ltvoff=-1.069952088e-08 wtvoff=2.849046863e-09 ptvoff=7.662282690e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.48 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.510960035e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.246677217e-08 wvth0=-1.352619098e-08 pvth0=-4.543245226e-14 k1=8.393317282e-01 lk1=-3.485796441e-07 wk1=-5.081662658e-07 pk1=6.873262002e-13 k2=-1.511863757e-01 lk2=1.186668036e-07 wk2=2.000365927e-07 pk2=-2.486705663e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.189402704e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.406838686e-07 wvoff=-1.558569208e-07 pvoff=-2.029185255e-13 nfactor=1.857754434e-01 lnfactor=1.020890666e-05 wnfactor=3.385652947e-06 pnfactor=-1.352824427e-11 eta0=0.08 etab=-0.07 u0=3.396287124e-02 lu0=1.193389280e-08 wu0=-5.209201394e-09 pu0=-2.154643820e-14 ua=-1.252734076e-09 lua=3.035089810e-15 wua=1.281001233e-15 pua=-6.132396179e-21 ub=2.217533366e-18 lub=-3.208534823e-24 wub=-1.627191798e-24 pub=6.937183691e-30 uc=2.395696424e-10 luc=-2.813594101e-16 wuc=-3.100019084e-16 puc=5.010287423e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=-2.078562241e-01 la0=5.272529140e-06 wa0=1.933469002e-06 pa0=-7.257488530e-12 ags=1.499051423e-01 lags=2.871477783e-06 wags=1.272072030e-07 pags=-3.165002513e-12 a1=0.0 a2=0.42385546 b0=-8.283076856e-24 lb0=3.264763146e-29 wb0=1.060757328e-29 pb0=-4.180960158e-35 b1=0.0 keta=-9.182995381e-02 lketa=2.336954727e-07 wketa=1.532262389e-07 pketa=-3.904318619e-13 dwg=0.0 dwb=0.0 pclm=3.647887870e-01 lpclm=-4.353553759e-08 wpclm=1.858726356e-07 ppclm=1.730079845e-13 pdiblc1=0.39 pdiblc2=4.380020132e-03 lpdiblc2=-1.741836728e-09 wpdiblc2=-3.752937327e-09 ppdiblc2=1.179663275e-14 pdiblcb=-0.025 drout=0.56 pscbe1=1.161900409e+09 lpscbe1=-7.681771935e+02 wpscbe1=-6.016933678e+02 ppscbe1=1.252128027e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.743289534e-01 lkt1=-7.883670925e-08 wkt1=1.007195875e-07 pkt1=1.109076414e-13 kt2=-1.008793767e-01 lkt2=-2.651400003e-08 wkt2=9.895336132e-08 pkt2=4.865244433e-14 at=1.526278299e+05 lat=-4.977241469e-02 wat=1.963153599e-02 pat=-7.737742426e-8 ute=-2.563567379e+00 lute=-4.986823275e-06 wute=1.068604993e-06 pute=9.635076550e-12 ua1=2.078181642e-09 lua1=-2.110888285e-14 wua1=-3.476694274e-15 pua1=3.759300911e-20 ub1=-3.596737599e-18 lub1=1.997524848e-23 wub1=5.614403551e-24 pub1=-3.434164863e-29 uc1=6.072844727e-11 luc1=4.137088959e-16 wuc1=-8.635020052e-17 puc1=-5.882875215e-22 kt1l=0.0 prt=0.0 tvoff=-3.218331638e-03 ltvoff=5.437299750e-09 wtvoff=7.598854993e-09 ptvoff=-1.105901956e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.49 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.753928194e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.529484421e-08 wvth0=-5.012265952e-08 pvth0=2.561907906e-14 k1=7.257372875e-01 lk1=-1.280376279e-07 wk1=-1.660725938e-07 pk1=2.315612530e-14 k2=-1.341797807e-01 lk2=8.564873752e-08 wk2=1.029264296e-07 pk2=-6.013254427e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.121918065e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.255823434e-07 wvoff=-3.880213034e-07 pvoff=2.478253731e-13 nfactor=7.204963244e+00 lnfactor=-3.418748186e-06 wnfactor=-5.294105261e-06 pnfactor=3.323384771e-12 eta0=1.529358871e-01 leta0=-1.416040037e-07 weta0=-2.441008415e-13 peta0=4.739183666e-19 etab=-5.646613875e-02 letab=-2.627580214e-8 u0=5.381567777e-02 lu0=-2.661005314e-08 wu0=-3.143546677e-08 pu0=2.937148885e-14 ua=2.246900721e-09 lua=-3.759402154e-15 wua=-4.076484055e-15 pua=4.269086502e-21 ub=-1.442301138e-18 lub=3.896982628e-24 wub=4.373473188e-24 pub=-4.713023371e-30 uc=9.969042798e-11 luc=-9.785873608e-18 wuc=-7.774368319e-17 puc=5.010264970e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.255379076e+05 lvsat=-8.841120999e-02 wvsat=-7.037427262e-02 pvsat=1.366306651e-7 a0=3.656203033e+00 la0=-2.229487810e-06 wa0=-2.937066941e-06 pa0=2.198588816e-12 ags=5.449709572e-01 lags=2.104463034e-06 wags=-2.508392541e-07 pags=-2.431030609e-12 a1=0.0 a2=0.42385546 b0=1.656615371e-23 lb0=-1.559680179e-29 wb0=-2.121514656e-29 pb0=1.997376347e-35 b1=0.0 keta=2.784170064e-01 lketa=-4.851338170e-07 wketa=-3.900384457e-07 pketa=6.643089175e-13 dwg=0.0 dwb=0.0 pclm=-7.492452152e-01 lpclm=2.119345881e-06 wpclm=1.514723106e-06 ppclm=-2.406936600e-12 pdiblc1=-6.362314151e-01 lpdiblc1=1.992413925e-06 wpdiblc1=1.376071480e-06 ppdiblc1=-2.671623514e-12 pdiblc2=1.092722770e-02 lpdiblc2=-1.445314856e-08 wpdiblc2=-7.824976357e-09 ppdiblc2=1.970243952e-14 pdiblcb=-1.895405684e-01 lpdiblcb=3.194532101e-07 wpdiblcb=2.401018180e-07 ppdiblcb=-4.661543183e-13 drout=1.236593378e+00 ldrout=-1.313596570e-06 wdrout=-6.702999833e-07 pdrout=1.301378033e-12 pscbe1=2.184201958e+09 lpscbe1=-2.752961339e+03 wpscbe1=-1.772653322e+03 ppscbe1=3.525530385e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.323601817e-08 lalpha0=2.198461440e-13 walpha0=1.464605049e-13 palpha0=-2.843510199e-19 alpha1=-4.317129657e-01 lalpha1=2.488427779e-06 walpha1=1.825874295e-06 palpha1=-3.544909381e-12 beta0=1.130964263e+01 lbeta0=4.951483130e-06 wbeta0=3.266069260e-06 pbeta0=-6.341027744e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-5.704107715e-01 lkt1=3.018533954e-07 wkt1=3.147039190e-07 pkt1=-3.045399423e-13 kt2=-1.897703609e-01 lkt2=1.460666012e-07 wkt2=2.426995743e-07 pkt2=-2.304288156e-13 at=2.424208118e+05 lat=-2.241042319e-01 wat=-1.373183800e-01 pat=2.273386404e-7 ute=-8.495401006e+00 lute=6.529748666e-06 wute=1.109120665e-05 pute=-9.823664251e-12 ua1=-1.972640126e-08 lua1=2.122440959e-14 wua1=3.273698888e-14 pua1=-3.271534974e-20 ub1=1.631254119e-17 lub1=-1.867833756e-23 wub1=-2.676781816e-23 pub1=2.852798146e-29 uc1=6.413391944e-10 luc1=-7.135387411e-16 wuc1=-9.182139546e-16 puc1=1.026764311e-21 kt1l=0.0 prt=0.0 tvoff=-1.658690061e-03 ltvoff=2.409277463e-09 wtvoff=3.687655584e-09 ptvoff=-3.465480663e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.50 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.012135010e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.014966085e-09 wvth0=-4.189671497e-08 pvth0=1.787446743e-14 k1=5.639451927e-01 lk1=2.428736434e-08 wk1=-2.036748725e-07 pk1=5.855814419e-14 k2=-3.320023220e-02 lk2=-9.422093717e-09 wk2=5.569364070e-08 pk2=-1.566353476e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.538418384e-01 ldsub=9.994642293e-08 wdsub=7.561656833e-08 pdsub=-7.119194045e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.075034106e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.390537411e-08 wvoff=-1.501690090e-08 pvoff=-1.033530498e-13 nfactor=1.031687874e+00 lnfactor=2.393304149e-06 wnfactor=8.269085289e-07 pnfactor=-2.439464018e-12 eta0=-4.278902942e-01 leta0=4.052357144e-07 weta0=4.882016829e-13 peta0=-2.155342084e-19 etab=-1.574825641e-01 letab=6.882974807e-08 wetab=-1.430811294e-09 petab=1.347088802e-15 u0=2.840727283e-02 lu0=-2.688395608e-09 wu0=-2.581985614e-10 pu0=1.852732054e-17 ua=-1.589862290e-09 lua=-1.471434945e-16 wua=3.614567046e-16 pua=9.082740857e-23 ub=2.673258171e-18 lub=2.224115675e-26 wub=-4.750923081e-25 pub=-1.481668361e-31 uc=1.058799697e-10 luc=-1.561324046e-17 wuc=-5.412774353e-17 puc=2.786857313e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.208725725e+04 lvsat=8.823525592e-02 wvsat=1.706147279e-01 pvsat=-9.025710506e-8 a0=1.101094316e+00 la0=1.761112748e-07 wa0=-1.133237181e-06 pa0=5.003083499e-13 ags=3.949146732e+00 lags=-1.100520799e-06 wags=-4.925973735e-06 pags=1.970543053e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.040468365e-01 lketa=1.573963365e-07 wketa=5.762211604e-07 pketa=-2.454109740e-13 dwg=0.0 dwb=0.0 pclm=2.743924296e+00 lpclm=-1.169424309e-06 wpclm=-2.419551617e-06 ppclm=1.297127972e-12 pdiblc1=1.381816268e+00 lpdiblc1=9.245028424e-08 wpdiblc1=-1.113550625e-06 ppdiblc1=-3.276791570e-13 pdiblc2=-7.917222451e-03 lpdiblc2=3.288637436e-09 wpdiblc2=2.232544433e-08 ppdiblc2=-8.683759449e-15 pdiblcb=3.040811369e-01 lpdiblcb=-1.452847148e-07 wpdiblcb=-4.802036361e-07 ppdiblcb=2.120031825e-13 drout=-1.181694435e+00 ldrout=9.631875495e-07 wdrout=1.340599967e-06 pdrout=-5.918561169e-13 pscbe1=-2.099509148e+09 lpscbe1=1.280092696e+03 wpscbe1=3.713204199e+03 ppscbe1=-1.639327669e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.122012203e-05 lalpha0=1.070506841e-11 walpha0=1.440437260e-11 palpha0=-1.370797565e-17 alpha1=3.413425931e+00 lalpha1=-1.131716661e-06 walpha1=-3.651748590e-06 palpha1=1.612195878e-12 beta0=4.094771402e+00 lbeta0=1.174418338e-05 wbeta0=1.250566423e-05 pbeta0=-1.503997705e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.011770546e-01 lkt1=-4.577497985e-08 wkt1=-5.505844492e-08 pkt1=4.358614663e-14 kt2=-3.105617084e-02 lkt2=-3.360586677e-09 wkt2=-6.482159624e-09 pkt2=4.172298272e-15 at=-2.335534459e+04 lat=2.612029843e-02 wat=1.799167076e-01 pat=-7.133375334e-8 ute=-1.757711648e+00 lute=1.863084626e-07 wute=1.112986939e-06 pute=-4.293100885e-13 ua1=4.524628971e-09 lua1=-1.607595861e-15 wua1=-4.025681542e-15 pua1=1.896189786e-21 ub1=-6.400284481e-18 lub1=2.705469831e-24 wub1=7.113757519e-24 pub1=-3.371047697e-30 uc1=-2.999409901e-10 luc1=1.726633747e-16 wuc1=3.833040672e-16 puc1=-1.985966853e-22 kt1l=0.0 prt=0.0 tvoff=-1.562006794e-04 ltvoff=9.947047457e-10 wtvoff=8.873027468e-10 ptvoff=-8.289876719e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.51 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.405887168e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.775002741e-08 wvth0=1.301831132e-07 pvth0=-5.809636760e-14 k1=7.957891642e-01 lk1=-7.806850328e-08 wk1=-6.345118851e-07 pk1=2.487666536e-13 k2=-1.403780741e-01 lk2=3.789542301e-08 wk2=2.206578426e-07 pk2=-8.849292039e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-3.601203002e-02 ldsub=1.837642479e-07 wdsub=3.049137622e-07 pdsub=-1.724234414e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-2.419113676e-03 lcdscd=3.452029220e-09 wcdscd=1.329743493e-08 pcdscd=-5.870631357e-15 cit=0.0 voff='-1.470582626e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.307108747e-08 wvoff=-1.995212868e-07 pvoff=-2.189694645e-14 nfactor=4.506873647e+00 lnfactor=8.590582831e-07 wnfactor=-1.571440256e-06 pnfactor=-1.380626606e-12 eta0=-6.527533278e-01 leta0=5.045095957e-07 weta0=1.943402877e-06 peta0=-8.579851627e-13 etab=-1.036035055e-01 letab=4.504289800e-08 wetab=1.751285417e-07 petab=-7.660139371e-14 u0=5.152080999e-02 lu0=-1.289269867e-08 wu0=-4.316623265e-08 pu0=1.896182366e-14 ua=3.477219062e-10 lua=-1.002559791e-15 wua=-2.657366670e-15 pua=1.423595665e-21 ub=2.195735225e-18 lub=2.330608520e-25 wub=-2.696374660e-25 pub=-2.388722725e-31 uc=1.099136038e-10 luc=-1.739403344e-17 wuc=-5.619167674e-17 puc=2.877977075e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.484487797e+05 lvsat=-4.713456880e-03 wvsat=-7.277957962e-02 pvsat=1.719807418e-8 a0=1.5 ags=5.430637904e+00 lags=-1.754578411e-06 wags=-5.703942656e-06 pags=2.314005440e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.543213828e-01 lketa=4.714604487e-08 wketa=2.076239100e-07 pketa=-8.268044826e-14 dwg=0.0 dwb=0.0 pclm=-2.714838865e-01 lpclm=1.618361877e-07 wpclm=1.244421652e-06 ppclm=-3.204649303e-13 pdiblc1=3.161737994e+00 lpdiblc1=-6.933602388e-07 wpdiblc1=-4.077768419e-06 ppdiblc1=9.809815003e-13 pdiblc2=1.079922882e-02 lpdiblc2=-4.974413768e-09 wpdiblc2=-1.844373716e-08 ppdiblc2=9.315263408e-15 pdiblcb=4.124239282e-01 lpdiblcb=-1.931165404e-07 wpdiblcb=-4.833793545e-07 ppdiblcb=2.134052177e-13 drout=-1.599597686e-01 ldrout=5.121059984e-07 wdrout=1.972664701e-06 pdrout=-8.709038483e-13 pscbe1=7.799614894e+08 lpscbe1=8.846721910e+00 wpscbe1=3.407813243e+01 ppscbe1=-1.504501837e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.282198546e-05 lalpha0=9.081454132e-14 walpha0=-1.637358642e-11 palpha0=-1.199376299e-19 alpha1=0.85 beta0=2.833111261e+01 lbeta0=1.044178050e-06 wbeta0=-1.898338038e-05 pbeta0=-1.138004704e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.371787784e-01 lkt1=1.426787721e-08 wkt1=5.582251428e-08 pkt1=-5.366244526e-15 kt2=-8.266258659e-02 lkt2=1.942292338e-08 wkt2=5.198056009e-08 pkt2=-2.163817400e-14 at=5.993417828e+04 lat=-1.065085986e-02 wat=8.445761554e-03 pat=4.368268758e-9 ute=-4.569275671e+00 lute=1.427574617e-06 wute=4.372894882e-06 pute=-1.868513807e-12 ua1=-5.903002580e-09 lua1=2.996057482e-15 wua1=1.005620064e-14 pua1=-4.320764051e-21 ub1=5.651304385e-18 lub1=-2.615137931e-24 wub1=-9.468718855e-24 pub1=3.949883468e-30 uc1=3.472775694e-10 luc1=-1.130745582e-16 wuc1=-5.004527604e-16 puc1=1.915695815e-22 kt1l=0.0 prt=0.0 tvoff=2.311535556e-04 ltvoff=8.236932739e-10 wtvoff=2.165696634e-09 ptvoff=-1.393380675e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.52 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.138420413e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.672637274e-08 wvth0=-5.183773770e-07 pvth0=6.609388644e-14 k1=-5.126107054e-01 lk1=1.724717542e-07 wk1=1.818093011e-06 pk1=-2.208728475e-13 k2=3.272797209e-01 lk2=-5.165449754e-08 wk2=-7.327830892e-07 pk2=9.407766987e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.730741775e+00 ldsub=-1.545443713e-07 wdsub=-1.629096067e-06 pdsub=1.979123648e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=3.913590781e-02 lcdscd=-4.505175625e-09 wcdscd=-4.749083903e-08 pcdscd=5.769472071e-15 cit=0.0 voff='1.545881989e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.468998684e-08 wvoff=-6.664336443e-07 pvoff=6.751023324e-14 nfactor=1.904442631e+01 lnfactor=-1.924679526e-06 wnfactor=-2.216850789e-05 pnfactor=2.563423486e-12 eta0=5.420459197e+00 leta0=-6.584255779e-07 weta0=-6.940724562e-06 peta0=8.432008642e-13 etab=4.364202597e-01 letab=-5.836409270e-08 wetab=-6.152389968e-07 petab=7.474292477e-14 u0=-1.008900091e-01 lu0=1.629183943e-08 wu0=1.769206434e-07 pu0=-2.318173189e-14 ua=-1.284335917e-08 lua=1.523347560e-15 wua=1.482481447e-14 pua=-1.923997273e-21 ub=6.901476871e-18 lub=-6.680227927e-25 wub=-5.508787724e-24 pub=7.643516538e-31 uc=2.905883578e-11 luc=-1.911477337e-18 wuc=1.069654640e-16 puc=-2.462537512e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.070567827e+04 lvsat=1.208811864e-02 wvsat=1.125178058e-01 pvsat=-1.828378096e-8 a0=1.5 ags=-1.237921116e+01 lags=1.655758347e-06 wags=1.745400395e-05 pags=-2.120417123e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.513665796e-01 lketa=-3.053752029e-08 wketa=-6.131910891e-07 pketa=7.449413265e-14 dwg=0.0 dwb=0.0 pclm=1.324694105e+00 lpclm=-1.438095512e-07 wpclm=-1.173937228e-06 ppclm=1.426169380e-13 pdiblc1=-1.875697085e+00 lpdiblc1=2.712380546e-07 wpdiblc1=2.859227667e-06 ppdiblc1=-3.473561324e-13 pdiblc2=-5.611053677e-02 lpdiblc2=7.837869604e-09 wpdiblc2=8.262208507e-08 ppdiblc2=-1.003742663e-14 pdiblcb=-1.451344888e+00 lpdiblcb=1.637690951e-07 wpdiblcb=1.726354838e-06 ppdiblcb=-2.097279438e-13 drout=6.004697136e+00 ldrout=-6.683394937e-07 wdrout=-7.045231076e-06 pdrout=8.558969424e-13 pscbe1=8.864570303e+08 lpscbe1=-1.154568324e+01 wpscbe1=-1.217076158e+02 ppscbe1=1.478577142e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.632000955e-05 lalpha0=-4.408728100e-12 walpha0=-4.650357428e-11 palpha0=5.649533225e-18 alpha1=0.85 beta0=6.859093906e+01 lbeta0=-6.665015078e-06 wbeta0=-6.845650031e-05 pbeta0=8.335405139e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.350500270e-01 lkt1=1.386025112e-08 wkt1=7.604264920e-08 pkt1=-9.238117280e-15 kt2=1.014654587e-01 lkt2=-1.583501950e-08 wkt2=-1.669232068e-07 pkt2=2.027883270e-14 at=-1.994215712e+05 lat=3.901213519e-02 wat=2.654953587e-01 pat=-4.485313041e-8 ute=1.018382254e+01 lute=-1.397437148e-06 wute=-1.473093796e-05 pute=1.789602729e-12 ua1=2.669446067e-08 lua1=-3.245900367e-15 wua1=-3.421632022e-14 pua1=4.156803878e-21 ub1=-2.312820516e-17 lub1=2.895735233e-24 wub1=3.052509098e-23 pub1=-3.708371203e-30 uc1=-9.208119192e-10 luc1=1.297468256e-16 wuc1=1.367712631e-15 puc1=-1.661579367e-22 kt1l=0.0 prt=0.0 tvoff=1.092886002e-02 ltvoff=-1.224767746e-09 wtvoff=-1.348185738e-08 ptvoff=1.602906852e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.53 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='3.422268371e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.566791574e-8 k1=0.90707349 k2=-9.790916945e-02 wk2=4.160795068e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-2.132730102e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.107298329e-7 nfactor=3.201617049e+00 wnfactor=-1.067940858e-6 eta0=0.00069413878 etab=-0.043998 u0=3.321465672e-02 wu0=-1.389749110e-8 ua=-3.040743130e-10 wua=-1.012378895e-15 ub=1.402713287e-18 wub=7.828973571e-25 uc=1.332469903e-11 wuc=8.669532994e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.602078319e+05 wvsat=-3.798332985e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=0.0 dwg=0.0 dwb=0.0 pclm=0.14094 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.372852629e+01 wbeta0=1.555631257e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=1.217029632e+05 wat=-1.037087504e-1 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=8.473053890e-04 wtvoff=-2.876880737e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.54 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='7.207531070e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.579205731e-06 wvth0=-2.266097733e-07 pvth0=4.518935621e-12 k1=4.897843500e-01 lk1=-3.244154722e-07 wk1=1.038770584e-07 pk1=-2.071462906e-12 k2=5.812723687e-03 lk2=-2.002040799e-07 wk2=-6.113878991e-08 pk2=1.219198323e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.835960858e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.825534760e-06 wvoff=-1.482108807e-07 pvoff=2.955545202e-12 nfactor=2.671654900e+00 lnfactor=3.943448818e-07 wnfactor=8.773490376e-08 pnfactor=-1.749564355e-12 eta0=0.08 etab=-0.07 u0=5.533900048e-02 lu0=-5.160039071e-07 wu0=-3.065069419e-08 pu0=6.112203890e-13 ua=1.015309237e-09 lua=-3.342018141e-14 wua=-2.212156907e-15 pua=4.411369599e-20 ub=3.777488064e-19 lub=2.253470064e-23 wub=1.567923842e-24 pub=-3.126673134e-29 uc=1.922537500e-10 luc=-3.319355067e-15 wuc=-1.408971056e-16 puc=2.809697660e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.319217779e+00 la0=3.729700146e-07 wa0=5.055590374e-08 pa0=-1.008159847e-12 ags=1.049379284e+00 lags=-1.399049360e-05 wags=-7.197779041e-07 pags=1.435344100e-11 a1=0.0 a2=0.42385546 b0=-3.537902388e-07 lb0=7.055103094e-12 wb0=4.530751011e-13 pb0=-9.034990785e-18 b1=-1.252975424e-07 lb1=2.498619187e-12 wb1=1.604600423e-13 pb1=-3.199811687e-18 keta=-1.213584887e-02 lketa=2.114294293e-07 wketa=6.979226811e-09 pketa=-1.391761537e-13 dwg=0.0 dwb=0.0 pclm=4.104129173e-01 lpclm=-6.518511177e-06 wpclm=-4.186154435e-07 ppclm=8.347814005e-12 pdiblc1=0.39 pdiblc2=9.657938736e-03 lpdiblc2=-1.297705370e-07 wpdiblc2=-9.434233052e-09 ppdiblc2=1.881326263e-13 pdiblcb=-1.477906972e+01 lpdiblcb=2.504754043e-04 wpdiblcb=1.561654031e-05 ppdiblcb=-3.114170199e-10 drout=0.56 pscbe1=3.589501872e+09 lpscbe1=-5.639428454e+04 wpscbe1=-3.570413546e+03 ppscbe1=7.119935175e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-4.692117897e-01 lkt1=3.524294510e-06 wkt1=1.881558852e-07 pkt1=-3.752107951e-12 kt2=-1.027635862e-01 lkt2=1.637733068e-06 wkt2=7.249736065e-08 pkt2=-1.445705102e-12 at=-3.164046903e+04 lat=3.422766010e+00 wat=2.198082771e-01 pat=-4.383303681e-6 ute=-5.225301030e+00 lute=7.852161581e-05 wute=4.238531607e-06 pute=-8.452261870e-11 ua1=-3.798811025e-09 lua1=1.027467323e-13 wua1=4.962140455e-15 pua1=-9.895245442e-20 ub1=4.113851003e-19 lub1=-2.698970652e-23 wub1=-9.063009278e-25 pub1=1.807298726e-29 uc1=-6.643260193e-11 luc1=8.380265700e-16 wuc1=1.171328792e-16 puc1=-2.335803670e-21 kt1l=0.0 prt=0.0 tvoff=-2.448240066e-03 ltvoff=9.880687381e-08 wtvoff=5.168634631e-09 ptvoff=-1.030702551e-13 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.55 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.5412677+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.47351598 k2=-0.0042268531 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32528737+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.69143 eta0=0.08 etab=-0.07 u0=0.0294631 ua=-6.6060305e-10 ub=1.50779e-18 uc=2.5799e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.337921 ags=0.347802 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.0015333577 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0031503727 pdiblcb=-2.2185512 drout=0.56 pscbe1=761513800.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.29248 kt2=-0.020636654 at=140000.0 ute=-1.2877 ua1=1.3536e-9 ub1=-9.4206e-19 uc1=-2.4408323e-11 kt1l=0.0 prt=0.0 tvoff=0.0025066 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.56 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.352432372e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.784318709e-8 k1=4.570235807e-01 lk1=1.309741580e-7 k2=5.544201942e-03 lk2=-7.759669682e-08 pk2=2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.307139784e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.309533435e-8 nfactor=2.644073046e+00 lnfactor=3.760845895e-7 eta0=0.08 etab=-0.07 u0=3.026006847e-02 lu0=-6.329113941e-9 ua=-6.244195286e-10 lua=-2.873509285e-16 ub=1.508341808e-18 lub=-4.382175824e-27 uc=2.621482677e-11 luc=-3.302282496e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.472040802e+00 la0=-1.065110528e-6 ags=3.449154527e-01 lags=2.292347475e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.266158166e-02 lketa=8.837463479e-08 wketa=-3.469446952e-24 pketa=2.081668171e-29 dwg=0.0 dwb=0.0 pclm=-3.595206022e-01 lpclm=3.518488096e-06 ppclm=1.332267630e-27 pdiblc1=0.39 pdiblc2=2.958945564e-03 lpdiblc2=1.520215920e-9 pdiblcb=-4.380014036e+00 lpdiblcb=1.716522685e-5 drout=0.56 pscbe1=7.775608705e+08 lpscbe1=-1.274375856e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912679931e-01 lkt1=-9.625136186e-9 kt2=-2.057583293e-02 lkt2=-4.830096796e-10 at=140000.0 ute=-1.486942117e+00 lute=1.582278485e-6 ua1=1.253190644e-09 lua1=7.973994938e-16 ub1=-9.359408430e-19 lub1=-4.859519977e-26 uc1=-3.044225720e-11 luc1=4.791840401e-17 kt1l=0.0 prt=0.0 tvoff=3.100483403e-03 ltvoff=-4.716316731e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.57 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.405338818e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.699018540e-8 k1=4.425227574e-01 lk1=1.881289500e-7 k2=5.015087822e-03 lk2=-7.551120093e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.406433988e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.223200618e-8 nfactor=2.829511464e+00 lnfactor=-3.548183393e-7 eta0=0.08 etab=-0.07 u0=2.989519107e-02 lu0=-4.890954778e-9 ua=-2.524457553e-10 lua=-1.753480349e-15 ub=9.469171404e-19 lub=2.208465292e-24 uc=-2.499826731e-12 luc=1.098761223e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.301920981e+00 la0=-3.945856366e-7 ags=2.492367247e-01 lags=4.000398419e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.781896867e-02 lketa=-7.117888762e-08 wketa=1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.099301200e-01 lpclm=9.156024676e-8 pdiblc1=0.39 pdiblc2=1.449484798e-03 lpdiblc2=7.469734397e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.920594498e+08 lpscbe1=2.095650671e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.956806083e-01 lkt1=7.767124987e-9 kt2=-2.361021482e-02 lkt2=1.147696406e-8 at=1.679573984e+05 lat=-1.101936944e-1 ute=-1.729131731e+00 lute=2.536865458e-6 ua1=-6.366453136e-10 lua1=8.246161464e-15 pua1=-3.308722450e-36 ub1=7.873505320e-19 lub1=-6.840924028e-24 pub1=3.081487911e-45 uc1=-6.699354411e-12 luc1=-4.566391495e-17 kt1l=0.0 prt=0.0 tvoff=2.715344074e-03 ltvoff=-3.198295456e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.58 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.362538165e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.529987224e-8 k1=5.960571032e-01 lk1=-1.099558329e-7 k2=-5.380819107e-02 lk2=3.869337152e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.817728603e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.206432023e-8 nfactor=3.070984661e+00 lnfactor=-8.236351706e-7 eta0=1.529356965e-01 leta0=-1.416036336e-7 etab=-5.646613875e-02 letab=-2.627580214e-8 u0=2.926883936e-02 lu0=-3.674901700e-9 ua=-9.362807507e-10 lua=-4.258242786e-16 ub=1.972788590e-18 lub=2.167502343e-25 uc=3.898314970e-11 luc=2.933750431e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.058514000e+04 lvsat=1.827881888e-2 a0=1.362751876e+00 la0=-5.126879678e-7 ags=3.490995015e-01 lags=2.061576588e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.615014926e-02 lketa=3.360139927e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=4.335482071e-01 lpclm=2.398546614e-7 pdiblc1=4.382938821e-01 lpdiblc1=-9.376189605e-8 pdiblc2=4.816981855e-03 lpdiblc2=9.317860066e-10 pdiblcb=-2.053594806e-03 lpdiblcb=-4.455012444e-8 drout=7.131799511e-01 ldrout=-2.973967305e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.112978320e-08 lalpha0=-2.193458266e-15 alpha1=9.940473580e-01 lalpha1=-2.796659289e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.246696694e-01 lkt1=6.404898136e-8 kt2=-2.548917326e-04 lkt2=-3.386706874e-8 at=1.351937707e+05 lat=-4.658356992e-2 ute=1.653279544e-01 lute=-1.141201499e-6 ua1=5.836749498e-09 lua1=-4.321843936e-15 ub1=-4.589496361e-18 lub1=3.598148939e-24 uc1=-7.566143859e-11 luc1=8.822500601e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=1.220869082e-03 ltvoff=-2.967931822e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.59 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.684978458e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.942570059e-9 k1=4.049027258e-01 lk1=7.001333729e-8 k2=1.028895181e-02 lk2=-2.165319114e-08 pk2=6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.128881283e-01 ldsub=4.435516763e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.192295746e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.200651935e-9 nfactor=1.677391346e+00 lnfactor=4.884134251e-7 eta0=-4.278899130e-01 leta0=4.052355461e-07 weta0=2.151057110e-22 peta0=-3.989863995e-29 etab=-1.585998337e-01 letab=6.988164183e-8 u0=2.820565476e-02 lu0=-2.673928282e-9 ua=-1.307613599e-09 lua=-7.621960020e-17 ub=2.302275478e-18 lub=-9.345705799e-26 uc=6.361353909e-11 luc=6.148337522e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.113971808e+04 lvsat=1.775669138e-2 a0=2.161896904e-01 la0=5.667842783e-7 ags=1.026289696e-01 lags=4.382062139e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.590378199e-02 lketa=-3.423636824e-08 wketa=-1.387778781e-23 pketa=-6.938893904e-30 dwg=0.0 dwb=0.0 pclm=8.545824573e-01 lpclm=-1.565431908e-7 pdiblc1=5.122841739e-01 lpdiblc1=-1.634227199e-7 pdiblc2=9.515923317e-03 lpdiblc2=-3.492201595e-9 pdiblcb=-7.089281039e-02 lpdiblcb=2.026103329e-8 drout=-1.348675822e-01 ldrout=5.010281494e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.774043360e-08 lalpha0=9.975669317e-16 alpha1=5.619052840e-01 lalpha1=1.271897838e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.441702368e-01 lkt1=-1.174010751e-8 kt2=-3.611785884e-02 lkt2=-1.025872893e-10 at=1.171352160e+05 lat=-2.958169351e-02 wat=1.164153218e-16 ute=-8.886197162e-01 lute=-1.489245227e-7 ua1=1.381117374e-09 lua1=-1.269286706e-16 ub1=-8.454041415e-19 lub1=7.313853160e-26 uc1=-6.324712557e-13 luc1=1.758628368e-17 kt1l=0.0 prt=0.0 tvoff=5.366624904e-04 ltvoff=3.473777448e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.60 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.422440817e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.761536061e-8 k1=3.003213912e-01 lk1=1.161845324e-7 k2=3.192579033e-02 lk2=-3.120555244e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.020842867e-01 ldsub=4.912491246e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380512e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-3.028573421e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.027459537e-9 nfactor=3.279791818e+00 lnfactor=-2.190239498e-7 eta0=8.647808876e-01 leta0=-1.654605150e-7 etab=3.314814661e-02 letab=-1.477240703e-08 wetab=-1.214306433e-23 petab=-5.746271514e-30 u0=1.781383355e-02 lu0=1.913915293e-9 ua=-1.727321252e-09 lua=1.090754525e-16 ub=1.985184914e-18 lub=4.653398671e-26 uc=6.603552112e-11 luc=5.079066363e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.161779340e+04 lvsat=8.715907823e-3 a0=1.5 ags=9.766318688e-01 lags=5.234616997e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=7.804747120e-03 lketa=-1.741617773e-08 pketa=6.938893904e-30 dwg=0.0 dwb=0.0 pclm=7.002407399e-01 lpclm=-8.840348330e-8 pdiblc1=-2.244639283e-02 lpdiblc1=7.265333909e-08 ppdiblc1=-2.775557562e-29 pdiblc2=-3.602829819e-03 lpdiblc2=2.299544252e-09 ppdiblc2=8.673617380e-31 pdiblcb=3.497017526e-02 lpdiblcb=-2.647599279e-08 ppdiblcb=-1.387778781e-29 drout=1.380423965e+00 ldrout=-1.679518545e-7 pscbe1=8.065718914e+08 lpscbe1=-2.901398061e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.643392960e-08 lalpha0=-2.840489843e-15 alpha1=0.85 beta0=1.350766576e+01 lbeta0=1.555506343e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.935889616e-01 lkt1=1.007756764e-8 kt2=-4.207281522e-02 lkt2=2.526442581e-9 at=6.652917321e+04 lat=-7.239834088e-3 ute=-1.154637522e+00 lute=-3.148138564e-8 ua1=1.949526982e-09 lua1=-3.778735547e-16 pua1=2.067951531e-37 ub1=-1.742481539e-18 lub1=4.691856435e-25 uc1=-4.350819919e-11 luc1=3.651531730e-17 puc1=-1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=1.922269063e-03 ltvoff=-2.643481584e-10 wtvoff=1.734723476e-24 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.61 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.150170992e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.248762530e-07 wvth0=-5.334255450e-07 pvth0=1.021435239e-13 k1=0.90707349 k2=-4.948307424e-01 lk2=6.966094899e-08 wk2=3.200378777e-07 pk2=-6.128277305e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586385734e-01 ldsub=-1.641693841e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-4.716902851e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.830168539e-08 wvoff=1.355986232e-07 pvoff=-2.596523796e-14 nfactor=-7.024897231e-01 lnfactor=5.435272134e-07 wnfactor=3.120024684e-06 pnfactor=-5.974410466e-13 eta0=6.941421173e-04 leta0=-4.054385601e-16 etab=-0.043998 u0=5.651529525e-02 lu0=-5.496872801e-09 wu0=-2.465762635e-08 pu0=4.721590240e-15 ua=-1.435491382e-09 lua=5.319411799e-17 wua=2.155339330e-16 pua=-4.127173070e-23 ub=4.127938494e-18 lub=-3.637733252e-25 wub=-1.956905725e-24 pub=3.747200497e-31 uc=3.112993757e-10 luc=-4.188552809e-17 wuc=-2.544808030e-16 puc=4.872951105e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.215520877e+05 lvsat=-1.616469046e-02 wvsat=-9.346725325e-02 pvsat=1.789767046e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.931507543e-01 lketa=7.850978741e-08 wketa=3.402616332e-07 pketa=-6.515533910e-14 dwg=0.0 dwb=0.0 pclm=3.311601613e-01 lpclm=-1.772971963e-08 wpclm=9.841413392e-08 ppclm=-1.884492885e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.020562730e-08 lalpha0=1.374977235e-14 walpha0=7.328712100e-14 palpha0=-1.403345765e-20 alpha1=0.85 beta0=1.670262989e+01 lbeta0=-4.562402672e-07 wbeta0=-2.006671170e-06 pbeta0=3.842494357e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-4.119265193e-01 lkt1=3.273755321e-08 wkt1=1.744931452e-07 pkt1=-3.341299441e-14 kt2=-0.028878939 at=1.441498091e+05 lat=-2.210309918e-02 wat=-1.744931452e-01 pat=3.341299441e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-2.228919154e-03 ltvoff=5.305462684e-10 wtvoff=3.368415676e-09 ptvoff=-6.450044441e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.62 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-6.128725966e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.930886042e-08 wvth0=1.248798814e-06 pvth0=-1.143717845e-13 k1=0.90707349 k2=4.705298602e-01 lk2=-4.761684918e-08 wk2=-6.863532607e-07 pk2=6.097966080e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-2.521352420e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.628821424e-09 wvoff=-6.096161519e-08 pvoff=-2.085920838e-15 nfactor=1.149277424e+01 lnfactor=-9.380266239e-07 wnfactor=-1.168586207e-05 pnfactor=1.201266911e-12 eta0=0.00069413878 etab=-0.043998 u0=-2.425311891e-02 lu0=4.315358761e-09 wu0=5.969758134e-08 pu0=-5.526386521e-15 ua=-8.219433528e-10 lua=-2.134337788e-17 wua=-3.491792306e-16 pua=2.733301270e-23 ub=-2.268167356e-18 lub=4.132639901e-25 wub=5.483944577e-24 pub=-5.292390902e-31 uc=-3.826463609e-10 luc=4.241916367e-17 wuc=5.937885404e-16 puc=-5.432333841e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.431768438e+04 lvsat=7.796528265e-03 wvsat=1.360419416e-01 pvsat=-9.984483585e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.199624958e-01 lketa=-5.671788889e-08 wketa=-7.939438109e-07 pketa=7.263474348e-14 dwg=0.0 dwb=0.0 pclm=1.852197268e-01 wpclm=-5.670603505e-8 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.635303837e-07 lalpha0=-1.221616068e-14 walpha0=-1.710032823e-13 palpha0=1.564440629e-20 alpha1=0.85 beta0=1.019381092e+01 lbeta0=3.344901139e-07 wbeta0=4.682232731e-06 pbeta0=-4.283587436e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=9.696874501e-02 lkt1=-2.908609687e-08 wkt1=-4.071506722e-07 pkt1=3.724858640e-14 kt2=-0.028878939 at=-2.772089980e+05 lat=2.908609687e-02 wat=4.071506722e-01 pat=-3.724858640e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=1.077251906e-02 ltvoff=-1.048946454e-09 wtvoff=-1.299823431e-08 ptvoff=1.343314396e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.63 nmos lmin=2.0e-05 lmax=0.0001 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.530635827e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.411773234e-06 wvth0=4.660272133e-08 pvth0=-4.657545222e-12 k1=7.182563689e-01 lk1=-1.501607324e-05 wk1=-1.293087952e-07 pk1=1.292331314e-11 k2=-1.076069596e-01 lk2=6.342897704e-06 wk2=5.462096828e-08 pk2=-5.458900736e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.325925897e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.482125537e-07 wvoff=3.859719141e-09 pvoff=-3.857460665e-13 nfactor=2.828652003e+00 lnfactor=-8.419270935e-06 wnfactor=-7.250136328e-08 pnfactor=7.245893984e-12 eta0=0.08 etab=-0.07 u0=2.084826226e-02 lu0=5.285643084e-07 wu0=4.551656935e-09 pu0=-4.548993579e-13 ua=-1.679669510e-09 lua=6.252493374e-14 wua=5.384246416e-16 pua=-5.381095878e-20 ub=2.349925937e-18 lub=-5.166934224e-23 wub=-4.449432476e-25 pub=4.446828935e-29 uc=8.469205205e-11 luc=-3.613389629e-15 wuc=-3.111619476e-17 puc=3.109798743e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.401841381e+00 la0=-3.921841967e-06 wa0=-3.377238853e-08 pa0=3.375262696e-12 ags=3.402338103e-01 lags=4.643471059e-07 wags=3.998659561e-09 pags=-3.996319785e-13 a1=0.0 a2=0.42385546 b0=1.868555482e-07 lb0=-1.146454253e-11 wb0=-9.872528976e-14 pb0=9.866752164e-18 b1=6.617633389e-08 lb1=-4.060256180e-12 wb1=-3.496432299e-14 pb1=3.494386396e-18 keta=-9.337871537e-03 lketa=4.788467972e-07 wketa=4.123521605e-09 pketa=-4.121108768e-13 dwg=0.0 dwb=0.0 pclm=-8.911282433e-02 lpclm=1.059258066e-05 wpclm=9.121651323e-08 ppclm=-9.116313880e-12 pdiblc1=0.39 pdiblc2=-2.522001665e-03 lpdiblc2=3.480291475e-07 wpdiblc2=2.997003880e-09 ppdiblc2=-2.995250213e-13 pdiblcb=3.462903853e+00 lpdiblcb=-3.485862941e-04 wpdiblcb=-3.001801669e-06 ppdiblcb=3.000045195e-10 drout=0.56 pscbe1=-6.280954511e+08 lpscbe1=8.525962708e+04 wpscbe1=7.342012443e+02 ppscbe1=-7.337716337e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.766805622e-01 lkt1=-9.693762308e-07 wkt1=-8.347646584e-09 pkt1=8.342762042e-13 kt2=-4.363979890e-02 lkt2=1.411360463e-06 wkt2=1.215373141e-08 pkt2=-1.214661978e-12 at=2.306525122e+05 lat=-5.561994767e+00 wat=-4.789633286e-02 pat=4.786830680e-6 ute=-8.414306329e-01 lute=-2.738090567e-05 wute=-2.357868043e-07 pute=2.356488360e-11 ua1=7.511493048e-10 lua1=3.696342808e-14 wua1=3.183053435e-16 pua1=-3.181190903e-20 ub1=2.297484320e-20 lub1=-5.920981800e-23 wub1=-5.098769903e-25 pub1=5.095786409e-29 uc1=1.264029705e-10 luc1=-9.253043350e-15 wuc1=-7.968127675e-17 puc1=7.963465204e-21 kt1l=0.0 prt=0.0 tvoff=2.733231280e-03 ltvoff=-1.390498692e-08 wtvoff=-1.197408322e-10 ptvoff=1.196707670e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.64 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='8.456720386e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.417422793e-06 wvth0=-3.106848089e-07 pvth0=2.467299060e-12 k1=-3.711162034e-01 lk1=6.707634659e-06 wk1=8.620586346e-07 pk1=-6.846026578e-12 k2=3.525518767e-01 lk2=-2.833353288e-06 wk2=-3.641397885e-07 pk2=2.891811033e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.000760686e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.002151969e-07 wvoff=-2.573146094e-08 pvoff=2.043460368e-13 nfactor=2.217858309e+00 lnfactor=3.760862952e-06 wnfactor=4.833424219e-07 pnfactor=-3.838457077e-12 eta0=0.08 etab=-0.07 u0=5.919407019e-02 lu0=-2.361080835e-07 wu0=-3.034437957e-08 pu0=2.409794655e-13 ua=2.856333133e-09 lua=-2.792969946e-14 wua=-3.589497610e-15 pua=2.850594502e-20 ub=-1.398535020e-18 lub=2.308053945e-23 wub=2.966288317e-24 pub=-2.355673714e-29 uc=-1.774488880e-10 luc=1.614090257e-15 wuc=2.074412984e-16 puc=-1.647392167e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.117323119e+00 la0=1.751874987e-06 wa0=2.251492569e-07 pa0=-1.788019671e-12 ags=3.739208464e-01 lags=-2.074224527e-07 wags=-2.665773040e-08 pags=2.117019928e-13 a1=0.0 a2=0.42385546 b0=-6.448637691e-07 lb0=5.121176594e-12 wb0=6.581685984e-13 pb0=-5.226836710e-18 b1=-2.283834787e-07 lb1=1.813704198e-12 wb1=2.330954866e-13 pb1=-1.851124543e-18 keta=2.540107512e-02 lketa=-2.138994211e-07 wketa=-2.749014404e-08 pketa=2.183125940e-13 dwg=0.0 dwb=0.0 pclm=6.793481880e-01 lpclm=-4.731673857e-06 wpclm=-6.081100882e-07 ppclm=4.829297752e-12 pdiblc1=0.39 pdiblc2=2.272650383e-02 lpdiblc2=-1.554635713e-07 wpdiblc2=-1.998002587e-08 ppdiblc2=1.586710957e-13 pdiblcb=-2.182602101e+01 lpdiblcb=1.557124470e-04 wpdiblcb=2.001201113e-05 ppdiblcb=-1.589251062e-10 drout=0.56 pscbe1=5.557243271e+09 lpscbe1=-3.808521846e+04 wpscbe1=-4.894674962e+03 ppscbe1=3.887099268e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.470059969e-01 lkt1=4.330174407e-07 wkt1=5.565097723e-08 pkt1=-4.419514565e-13 kt2=5.875031023e-02 lkt2=-6.304504650e-07 wkt2=-8.102487608e-08 pkt2=6.434579190e-13 at=-1.728540803e+05 lat=2.484526299e+00 wat=3.193088857e-01 pat=-2.535787046e-6 ute=-2.827835944e+00 lute=1.223096804e-05 wute=1.571912029e-06 pute=-1.248331737e-11 ua1=3.432738831e-09 lua1=-1.651145192e-14 wua1=-2.122035623e-15 pua1=1.685211620e-20 ub1=-4.272525766e-18 lub1=2.644884725e-23 wub1=3.399179935e-24 pub1=-2.699453987e-29 uc1=-5.448784941e-10 luc1=4.133306577e-15 wuc1=5.312085116e-16 puc1=-4.218584958e-21 kt1l=0.0 prt=0.0 tvoff=1.724464799e-03 ltvoff=6.211315748e-09 wtvoff=7.982722143e-10 ptvoff=-6.339467614e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.65 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.352432372e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.784318709e-8 k1=4.570235807e-01 lk1=1.309741580e-7 k2=5.544201942e-03 lk2=-7.759669682e-08 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.307139784e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.309533435e-8 nfactor=2.644073046e+00 lnfactor=3.760845895e-7 eta0=0.08 etab=-0.07 u0=3.026006847e-02 lu0=-6.329113941e-9 ua=-6.244195286e-10 lua=-2.873509285e-16 ub=1.508341808e-18 lub=-4.382175824e-27 uc=2.621482677e-11 luc=-3.302282496e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.472040802e+00 la0=-1.065110528e-06 wa0=-1.776356839e-21 ags=3.449154527e-01 lags=2.292347475e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.266158166e-02 lketa=8.837463479e-08 wketa=-3.469446952e-24 dwg=0.0 dwb=0.0 pclm=-3.595206022e-01 lpclm=3.518488096e-06 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=2.958945564e-03 lpdiblc2=1.520215920e-9 pdiblcb=-4.380014036e+00 lpdiblcb=1.716522685e-5 drout=0.56 pscbe1=7.775608705e+08 lpscbe1=-1.274375856e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912679931e-01 lkt1=-9.625136186e-9 kt2=-2.057583293e-02 lkt2=-4.830096796e-10 at=140000.0 ute=-1.486942117e+00 lute=1.582278485e-06 wute=-1.776356839e-21 ua1=1.253190644e-09 lua1=7.973994938e-16 ub1=-9.359408430e-19 lub1=-4.859519977e-26 uc1=-3.044225720e-11 luc1=4.791840401e-17 kt1l=0.0 prt=0.0 tvoff=3.100483403e-03 ltvoff=-4.716316731e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.66 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.405338818e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.699018540e-8 k1=4.425227574e-01 lk1=1.881289500e-7 k2=5.015087822e-03 lk2=-7.551120093e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.406433988e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.223200618e-8 nfactor=2.829511464e+00 lnfactor=-3.548183393e-7 eta0=0.08 etab=-0.07 u0=2.989519107e-02 lu0=-4.890954778e-9 ua=-2.524457553e-10 lua=-1.753480349e-15 ub=9.469171404e-19 lub=2.208465292e-24 uc=-2.499826731e-12 luc=1.098761223e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.301920981e+00 la0=-3.945856366e-7 ags=2.492367247e-01 lags=4.000398419e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.781896867e-02 lketa=-7.117888762e-8 dwg=0.0 dwb=0.0 pclm=5.099301200e-01 lpclm=9.156024676e-8 pdiblc1=0.39 pdiblc2=1.449484798e-03 lpdiblc2=7.469734397e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.920594498e+08 lpscbe1=2.095650671e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.956806083e-01 lkt1=7.767124987e-9 kt2=-2.361021482e-02 lkt2=1.147696406e-8 at=1.679573984e+05 lat=-1.101936944e-1 ute=-1.729131731e+00 lute=2.536865458e-6 ua1=-6.366453136e-10 lua1=8.246161464e-15 ub1=7.873505320e-19 lub1=-6.840924028e-24 uc1=-6.699354411e-12 luc1=-4.566391495e-17 kt1l=0.0 prt=0.0 tvoff=2.715344074e-03 ltvoff=-3.198295456e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.67 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.362538165e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.529987224e-8 k1=5.960571032e-01 lk1=-1.099558329e-7 k2=-5.380819107e-02 lk2=3.869337152e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.817728603e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.206432023e-8 nfactor=3.070984661e+00 lnfactor=-8.236351706e-7 eta0=1.529356965e-01 leta0=-1.416036336e-7 etab=-5.646613875e-02 letab=-2.627580214e-8 u0=2.926883936e-02 lu0=-3.674901700e-9 ua=-9.362807507e-10 lua=-4.258242786e-16 ub=1.972788590e-18 lub=2.167502343e-25 uc=3.898314970e-11 luc=2.933750431e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.058514000e+04 lvsat=1.827881888e-2 a0=1.362751876e+00 la0=-5.126879678e-7 ags=3.490995015e-01 lags=2.061576588e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.615014926e-02 lketa=3.360139927e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=4.335482071e-01 lpclm=2.398546614e-7 pdiblc1=4.382938821e-01 lpdiblc1=-9.376189605e-8 pdiblc2=4.816981855e-03 lpdiblc2=9.317860066e-10 pdiblcb=-2.053594806e-03 lpdiblcb=-4.455012444e-8 drout=7.131799511e-01 ldrout=-2.973967305e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.112978320e-08 lalpha0=-2.193458266e-15 alpha1=9.940473580e-01 lalpha1=-2.796659289e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.246696694e-01 lkt1=6.404898136e-8 kt2=-2.548917326e-04 lkt2=-3.386706874e-8 at=1.351937707e+05 lat=-4.658356992e-2 ute=1.653279544e-01 lute=-1.141201499e-6 ua1=5.836749498e-09 lua1=-4.321843936e-15 ub1=-4.589496361e-18 lub1=3.598148939e-24 pub1=3.081487911e-45 uc1=-7.566143859e-11 luc1=8.822500601e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=1.220869082e-03 ltvoff=-2.967931822e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.68 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.684978458e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.942570059e-9 k1=4.049027258e-01 lk1=7.001333729e-8 k2=1.028895181e-02 lk2=-2.165319114e-08 pk2=6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.128881283e-01 ldsub=4.435516763e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.192295746e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.200651935e-9 nfactor=1.677391346e+00 lnfactor=4.884134251e-7 eta0=-4.278899130e-01 leta0=4.052355461e-07 weta0=1.873501354e-22 peta0=1.006139616e-28 etab=-1.585998338e-01 letab=6.988164183e-8 u0=2.820565476e-02 lu0=-2.673928282e-9 ua=-1.307613599e-09 lua=-7.621960020e-17 ub=2.302275478e-18 lub=-9.345705799e-26 uc=6.361353909e-11 luc=6.148337522e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.113971808e+04 lvsat=1.775669138e-2 a0=2.161896904e-01 la0=5.667842783e-7 ags=1.026289696e-01 lags=4.382062139e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.590378199e-02 lketa=-3.423636824e-08 wketa=1.387778781e-23 pketa=6.938893904e-30 dwg=0.0 dwb=0.0 pclm=8.545824573e-01 lpclm=-1.565431908e-7 pdiblc1=5.122841739e-01 lpdiblc1=-1.634227199e-7 pdiblc2=9.515923317e-03 lpdiblc2=-3.492201595e-9 pdiblcb=-7.089281039e-02 lpdiblcb=2.026103329e-8 drout=-1.348675822e-01 ldrout=5.010281494e-07 pdrout=2.220446049e-28 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.774043360e-08 lalpha0=9.975669317e-16 alpha1=5.619052840e-01 lalpha1=1.271897838e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.441702368e-01 lkt1=-1.174010751e-8 kt2=-3.611785884e-02 lkt2=-1.025872893e-10 at=1.171352160e+05 lat=-2.958169351e-2 ute=-8.886197162e-01 lute=-1.489245227e-7 ua1=1.381117374e-09 lua1=-1.269286706e-16 wua1=-1.654361225e-30 ub1=-8.454041415e-19 lub1=7.313853160e-26 uc1=-6.324712557e-13 luc1=1.758628368e-17 kt1l=0.0 prt=0.0 tvoff=5.366624904e-04 ltvoff=3.473777448e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.69 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.422440817e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.761536061e-8 k1=3.003213912e-01 lk1=1.161845324e-7 k2=3.192579033e-02 lk2=-3.120555244e-08 pk2=-1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.020842867e-01 ldsub=4.912491246e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380512e-03 lcdscd=-1.132138095e-09 wcdscd=-6.938893904e-24 cit=0.0 voff='-3.028573421e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.027459537e-9 nfactor=3.279791818e+00 lnfactor=-2.190239498e-07 wnfactor=3.552713679e-21 eta0=8.647808876e-01 leta0=-1.654605150e-7 etab=3.314814661e-02 letab=-1.477240703e-08 wetab=-7.806255642e-24 petab=-4.228388473e-30 u0=1.781383355e-02 lu0=1.913915293e-9 ua=-1.727321252e-09 lua=1.090754525e-16 ub=1.985184914e-18 lub=4.653398671e-26 uc=6.603552112e-11 luc=5.079066363e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.161779340e+04 lvsat=8.715907823e-3 a0=1.5 ags=9.766318688e-01 lags=5.234616997e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=7.804747120e-03 lketa=-1.741617773e-8 dwg=0.0 dwb=0.0 pclm=7.002407399e-01 lpclm=-8.840348330e-8 pdiblc1=-2.244639283e-02 lpdiblc1=7.265333909e-8 pdiblc2=-3.602829819e-03 lpdiblc2=2.299544252e-9 pdiblcb=3.497017526e-02 lpdiblcb=-2.647599279e-08 ppdiblcb=-6.938893904e-30 drout=1.380423965e+00 ldrout=-1.679518545e-7 pscbe1=8.065718914e+08 lpscbe1=-2.901398061e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.643392960e-08 lalpha0=-2.840489843e-15 alpha1=0.85 beta0=1.350766576e+01 lbeta0=1.555506343e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.935889616e-01 lkt1=1.007756764e-8 kt2=-4.207281522e-02 lkt2=2.526442581e-9 at=6.652917321e+04 lat=-7.239834088e-3 ute=-1.154637522e+00 lute=-3.148138564e-8 ua1=1.949526982e-09 lua1=-3.778735547e-16 ub1=-1.742481539e-18 lub1=4.691856435e-25 uc1=-4.350819919e-11 luc1=3.651531730e-17 kt1l=0.0 prt=0.0 tvoff=1.922269063e-03 ltvoff=-2.643481584e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.70 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.275286050e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.479755284e-8 k1=0.90707349 k2=-1.812624066e-01 lk2=9.617002643e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586385734e-01 ldsub=-1.641693841e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-3.388327780e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.861332788e-9 nfactor=2.354463893e+00 lnfactor=-4.183660682e-8 eta0=6.941421173e-04 leta0=-4.054385601e-16 etab=-0.043998 u0=3.235612098e-02 lu0=-8.707291566e-10 ua=-1.224314451e-09 lua=1.275669227e-17 ub=2.210591472e-18 lub=3.371786582e-27 uc=6.196288314e-11 luc=5.858919519e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.299742681e+05 lvsat=1.371179917e-3 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.597674847e-01 lketa=1.467155864e-8 dwg=0.0 dwb=0.0 pclm=4.275848609e-01 lpclm=-3.619369965e-08 wpclm=4.440892099e-22 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.16e-8 alpha1=0.85 beta0=1.473652343e+01 lbeta0=-7.975840524e-8 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.24096074 kt2=-0.028878939 at=-2.681597014e+04 lat=1.063445403e-2 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=1.071404250e-03 ltvoff=-1.014194588e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.71 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.062807568e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.852676324e-08 wvth0=5.148078884e-07 pvth0=-6.254195113e-14 k1=0.90707349 k2=-1.747193634e-01 lk2=8.822114501e-09 wk2=-2.779125511e-08 pk2=3.376248419e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587060922e-01 ldsub=-9.844282633e-12 wdsub=-8.270409654e-11 pdsub=1.004738987e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-8.697545346e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.773580614e-08 wvoff=-2.295289805e-07 pvoff=2.788455772e-14 nfactor=-8.199674913e+00 lnfactor=1.240343500e-06 wnfactor=8.412881691e-06 pnfactor=-1.022047345e-12 eta0=-1.069201800e-02 leta0=1.383258773e-09 weta0=1.162107706e-08 peta0=-1.411798168e-15 etab=-0.043998 u0=2.198606496e-02 lu0=3.890874693e-10 wu0=1.250439063e-08 pu0=-1.519108400e-15 ua=-2.111517827e-09 lua=1.205394816e-16 wua=9.670017442e-16 pua=-1.174771739e-22 ub=6.288043207e-18 lub=-4.919815149e-25 wub=-3.248797723e-24 pub=3.946834401e-31 uc=1.332303798e-10 luc=-2.799083581e-18 wuc=6.726823075e-17 puc=-8.172148281e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.507857807e+05 lvsat=-1.157127505e-03 wvsat=6.964555498e-03 pvsat=-8.460959892e-10 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=9.360371878e-06 lb0=-1.137154138e-12 wb0=-9.553495071e-12 pb0=1.160615902e-18 b1=-1.337704485e-08 lb1=1.625123670e-15 wb1=1.365304003e-14 pb1=-1.658653222e-21 keta=-6.008205577e-01 lketa=6.825333228e-08 wketa=4.520264386e-07 pketa=-5.491488392e-14 dwg=0.0 dwb=0.0 pclm=1.037428060e-01 lpclm=3.148576227e-09 wpclm=2.645191752e-08 ppclm=-3.213537651e-15 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.016080000e-09 lalpha0=3.111995095e-15 alpha1=0.85 beta0=1.806205013e+01 lbeta0=-4.837633423e-07 wbeta0=-3.348343989e-06 pbeta0=4.067769179e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-6.300171531e-01 lkt1=4.726490741e-08 wkt1=3.348343989e-07 pkt1=-4.067769179e-14 kt2=-0.028878939 at=3.349538889e+05 lat=-3.331551906e-02 wat=-2.176423593e-01 pat=2.644049966e-8 ute=-4.988788338e-01 lute=-9.963848819e-08 wute=-8.370859974e-07 pute=1.016942295e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-9.215998463e-03 ltvoff=1.148355947e-09 wtvoff=7.402686309e-09 ptvoff=-8.993227490e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.72 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.73 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.846759231e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.494228043e-7 k1=6.305414559e-01 lk1=-1.247015618e-6 k2=-7.055554732e-02 lk2=5.267483965e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.299744003e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.722198512e-8 nfactor=2.779471661e+00 lnfactor=-6.991816158e-7 eta0=0.08 etab=-0.07 u0=2.393581862e-02 lu0=4.389482771e-8 ua=-1.314436267e-09 lua=5.192407340e-15 ub=2.048104563e-18 lub=-4.290900539e-24 uc=6.358479239e-11 luc=-3.000753413e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.378932328e+00 la0=-3.256908852e-7 ags=3.429462482e-01 lags=3.856188526e-8 a1=0.0 a2=0.42385546 b0=1.198865520e-07 lb0=-9.520773746e-13 b1=4.245874728e-08 lb1=-3.371855471e-13 keta=-6.540735128e-03 lketa=3.976601774e-8 dwg=0.0 dwb=0.0 pclm=-2.723730757e-02 lpclm=8.796649638e-7 pdiblc1=0.39 pdiblc2=-4.890236744e-04 lpdiblc2=2.890221536e-8 pdiblcb=1.426671345e+00 lpdiblcb=-2.894848381e-05 wpdiblcb=-7.771561172e-22 ppdiblcb=-6.661338148e-27 drout=0.56 pscbe1=-1.300597360e+08 lpscbe1=7.080418754e+03 ppscbe1=-3.814697266e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.823430780e-01 lkt1=-8.050222454e-8 kt2=-3.539547575e-02 lkt2=1.172069763e-7 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.001373497e+00 lute=-2.273857916e-6 ua1=9.670675297e-10 lua1=3.069642201e-15 ub1=-3.228934776e-19 lub1=-4.917102269e-24 uc1=7.235222898e-11 luc1=-7.684225689e-16 wuc1=-5.169878828e-32 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=2.652006669e-03 ltvoff=-1.154745024e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.74 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.352432372e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.784318709e-8 k1=4.570235807e-01 lk1=1.309741580e-7 k2=5.544201942e-03 lk2=-7.759669682e-08 pk2=5.551115123e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.307139784e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.309533435e-8 nfactor=2.644073046e+00 lnfactor=3.760845895e-7 eta0=0.08 etab=-0.07 u0=3.026006847e-02 lu0=-6.329113941e-9 ua=-6.244195286e-10 lua=-2.873509285e-16 ub=1.508341808e-18 lub=-4.382175824e-27 uc=2.621482677e-11 luc=-3.302282496e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.472040802e+00 la0=-1.065110528e-6 ags=3.449154527e-01 lags=2.292347475e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.266158166e-02 lketa=8.837463479e-08 wketa=3.469446952e-24 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=-3.595206022e-01 lpclm=3.518488096e-06 wpclm=-2.220446049e-22 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=2.958945564e-03 lpdiblc2=1.520215920e-9 pdiblcb=-4.380014036e+00 lpdiblcb=1.716522685e-5 drout=0.56 pscbe1=7.775608705e+08 lpscbe1=-1.274375856e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912679931e-01 lkt1=-9.625136186e-9 kt2=-2.057583293e-02 lkt2=-4.830096796e-10 at=140000.0 ute=-1.486942117e+00 lute=1.582278485e-6 ua1=1.253190644e-09 lua1=7.973994938e-16 ub1=-9.359408430e-19 lub1=-4.859519977e-26 uc1=-3.044225720e-11 luc1=4.791840401e-17 kt1l=0.0 prt=0.0 tvoff=3.100483403e-03 ltvoff=-4.716316731e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.75 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.405338818e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.699018540e-8 k1=4.425227574e-01 lk1=1.881289500e-7 k2=5.015087822e-03 lk2=-7.551120093e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.406433988e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.223200618e-8 nfactor=2.829511464e+00 lnfactor=-3.548183393e-7 eta0=0.08 etab=-0.07 u0=2.989519107e-02 lu0=-4.890954778e-9 ua=-2.524457553e-10 lua=-1.753480349e-15 ub=9.469171404e-19 lub=2.208465292e-24 uc=-2.499826731e-12 luc=1.098761223e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.301920981e+00 la0=-3.945856366e-7 ags=2.492367247e-01 lags=4.000398419e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.781896867e-02 lketa=-7.117888762e-08 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=5.099301200e-01 lpclm=9.156024676e-8 pdiblc1=0.39 pdiblc2=1.449484798e-03 lpdiblc2=7.469734397e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.920594498e+08 lpscbe1=2.095650671e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.956806083e-01 lkt1=7.767124987e-9 kt2=-2.361021482e-02 lkt2=1.147696406e-8 at=1.679573984e+05 lat=-1.101936944e-01 wat=-2.328306437e-16 ute=-1.729131731e+00 lute=2.536865458e-6 ua1=-6.366453136e-10 lua1=8.246161464e-15 ub1=7.873505320e-19 lub1=-6.840924028e-24 pub1=-3.081487911e-45 uc1=-6.699354411e-12 luc1=-4.566391495e-17 kt1l=0.0 prt=0.0 tvoff=2.715344074e-03 ltvoff=-3.198295456e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.76 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.362538165e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.529987224e-8 k1=5.960571032e-01 lk1=-1.099558329e-7 k2=-5.380819107e-02 lk2=3.869337152e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.817728603e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.206432023e-8 nfactor=3.070984661e+00 lnfactor=-8.236351706e-7 eta0=1.529356965e-01 leta0=-1.416036336e-7 etab=-5.646613875e-02 letab=-2.627580214e-8 u0=2.926883936e-02 lu0=-3.674901700e-9 ua=-9.362807507e-10 lua=-4.258242786e-16 ub=1.972788590e-18 lub=2.167502343e-25 uc=3.898314970e-11 luc=2.933750431e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.058514000e+04 lvsat=1.827881888e-2 a0=1.362751876e+00 la0=-5.126879678e-7 ags=3.490995015e-01 lags=2.061576588e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.615014926e-02 lketa=3.360139927e-8 dwg=0.0 dwb=0.0 pclm=4.335482071e-01 lpclm=2.398546614e-7 pdiblc1=4.382938821e-01 lpdiblc1=-9.376189605e-8 pdiblc2=4.816981855e-03 lpdiblc2=9.317860066e-10 pdiblcb=-2.053594806e-03 lpdiblcb=-4.455012444e-8 drout=7.131799511e-01 ldrout=-2.973967305e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.112978320e-08 lalpha0=-2.193458266e-15 alpha1=9.940473580e-01 lalpha1=-2.796659289e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.246696694e-01 lkt1=6.404898136e-08 wkt1=-4.440892099e-22 kt2=-2.548917326e-04 lkt2=-3.386706874e-8 at=1.351937707e+05 lat=-4.658356992e-2 ute=1.653279544e-01 lute=-1.141201499e-6 ua1=5.836749498e-09 lua1=-4.321843936e-15 ub1=-4.589496361e-18 lub1=3.598148939e-24 wub1=6.162975822e-39 uc1=-7.566143859e-11 luc1=8.822500601e-17 wuc1=5.169878828e-32 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=1.220869082e-03 ltvoff=-2.967931822e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.77 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='7.561677608e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.689831969e-07 wvth0=4.241892208e-07 pvth0=-3.993682127e-13 k1=-1.895070522e-01 lk1=6.296418215e-07 wk1=5.115680760e-07 pk1=-4.816341816e-13 k2=1.797896551e-01 lk2=-1.812357303e-07 wk2=-1.458777293e-07 pk2=1.373418398e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.924112721e-01 ldsub=6.363384111e-08 wdsub=1.762303774e-08 pdsub=-1.659184331e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='8.113930453e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.061264716e-06 wvoff=-9.730500067e-07 pvoff=9.161129586e-13 nfactor=1.596653823e+01 lnfactor=-1.296461832e-05 wnfactor=-1.229769706e-05 pnfactor=1.157810962e-11 eta0=-4.278899128e-01 leta0=4.052355460e-07 weta0=-1.160077451e-16 peta0=1.092194772e-22 etab=-1.606986361e-01 letab=7.185763485e-08 wetab=1.806296458e-09 petab=-1.700602827e-15 u0=4.357291779e-02 lu0=-1.714199129e-08 wu0=-1.322555832e-08 pu0=1.245167800e-14 ua=-1.096653404e-09 lua=-2.748356712e-16 wua=-1.815590953e-16 pua=1.709353464e-22 ub=2.686925170e-18 lub=-4.555993582e-25 wub=-3.310418340e-25 pub=3.116712521e-31 uc=-1.043107990e-10 luc=1.642467509e-16 wuc=1.445210590e-16 puc=-1.360645537e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.433556872e+05 lvsat=-1.443822325e-01 wvsat=-1.482145739e-01 pvsat=1.395419464e-7 a0=-5.588560472e-01 la0=1.296478990e-06 wa0=6.670291633e-07 pa0=-6.279986188e-13 ags=-6.203516576e+00 lags=6.375353959e-06 wags=5.427270653e-06 pags=-5.109699338e-12 a1=0.0 a2=0.42385546 b0=4.892557602e-16 lb0=-4.606274487e-22 wb0=-4.210691634e-22 pb0=3.964307224e-28 b1=-2.408618580e-17 lb1=2.267680672e-23 wb1=2.072934226e-23 pb1=-1.951638552e-29 keta=2.106576318e-01 lketa=-1.893498113e-07 wketa=-1.417924353e-07 pketa=1.334955927e-13 dwg=0.0 dwb=0.0 pclm=5.309303398e-01 lpclm=1.481707468e-07 wpclm=2.785453692e-07 ppclm=-2.622465655e-13 pdiblc1=-2.203641250e-01 lpdiblc1=5.263553964e-07 wpdiblc1=6.305405707e-07 ppdiblc1=-5.936451198e-13 pdiblc2=-9.571235793e-04 lpdiblc2=6.368025435e-09 wpdiblc2=9.013439296e-09 ppdiblc2=-8.486026909e-15 pdiblcb=-5.383730653e-01 lpdiblcb=4.603871486e-07 wpdiblcb=4.023284668e-07 ppdiblcb=-3.787866189e-13 drout=-1.348682540e-01 ldrout=5.010287819e-07 wdrout=5.782008330e-13 pdrout=-5.443679889e-19 pscbe1=-1.638324720e+09 lpscbe1=2.295648587e+03 wpscbe1=2.098500280e+03 ppscbe1=-1.975708635e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.601930898e-05 lalpha0=-2.446970034e-11 walpha0=-2.236917562e-11 palpha0=2.106026568e-17 alpha1=5.619052840e-01 lalpha1=1.271897838e-7 beta0=4.178582480e+01 lbeta0=-2.629177309e-05 wbeta0=-2.403385845e-05 pbeta0=2.262754125e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.841628505e+00 lkt1=2.433730488e-06 wkt1=2.235455705e-06 pkt1=-2.104650250e-12 kt2=-3.859191364e-02 lkt2=2.226700666e-09 wkt2=2.129250729e-09 pkt2=-2.004659751e-15 at=-1.479863587e+05 lat=2.200265574e-01 wat=2.281721111e-01 pat=-2.148208482e-7 ute=-1.455018307e+00 lute=3.843318212e-07 wute=4.874607522e-07 pute=-4.589374737e-13 ua1=-3.781459853e-10 lua1=1.529393153e-15 wua1=1.514078344e-15 pua1=-1.425483564e-21 ub1=-5.239636594e-19 lub1=-2.294931821e-25 wub1=-2.766419650e-25 pub1=2.604545370e-31 uc1=-2.253648137e-10 luc1=2.291686378e-16 wuc1=1.934118454e-16 puc1=-1.820945446e-22 kt1l=0.0 prt=0.0 tvoff=-8.352185306e-03 ltvoff=8.716103501e-09 wtvoff=7.650026856e-09 ptvoff=-7.202393185e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.78 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.356857649e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.666671115e-08 wvth0=-6.150193037e-07 pvth0=5.942780192e-14 k1=1.489140946e+00 lk1=-1.114577688e-07 wk1=-1.023136151e-06 pk1=1.959162489e-13 k2=-3.314376233e-01 lk2=4.446395595e-08 wk2=3.127221814e-07 pk2=-6.512360034e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.430379993e-01 ldsub=4.128284982e-08 wdsub=-3.524607558e-08 pdsub=6.749130055e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380505e-03 lcdscd=-1.132138092e-09 wcdscd=6.154451948e-18 pcdscd=-2.717104319e-24 cit=0.0 voff='-1.716941717e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.495968461e-08 wvoff=1.217006263e-06 pvoff=-5.076622384e-14 nfactor=-1.314881340e+01 lnfactor=-1.105981878e-07 wnfactor=1.413898337e-05 pnfactor=-9.331468036e-14 eta0=8.647808877e-01 leta0=-1.654605150e-07 weta0=-3.877609345e-17 peta0=7.512279687e-23 etab=3.734575126e-02 letab=-1.557618955e-08 wetab=-3.612592886e-09 petab=6.917609541e-16 u0=-2.418717612e-03 lu0=3.162671860e-09 wu0=1.741278098e-08 pu0=-1.074719861e-15 ua=-2.292707264e-09 lua=2.532053636e-16 wua=4.865892945e-16 pua=-1.240428136e-22 ub=1.343125702e-18 lub=1.376692938e-25 wub=5.525767038e-25 pub=-7.843396165e-32 uc=4.018841974e-10 luc=-5.923125330e-17 wuc=-2.890421180e-16 puc=5.534751903e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-2.335067304e+05 lvsat=6.614584877e-02 wvsat=2.798125691e-01 pvsat=-4.942604494e-8 a0=3.050091473e+00 la0=-2.968208152e-07 wa0=-1.334058324e-06 pa0=2.554534918e-13 ags=1.358892296e+01 lags=-2.362731002e-06 wags=-1.085454131e-05 pags=2.078492696e-12 a1=0.0 a2=0.42385546 b0=-9.785115205e-16 lb0=1.873712570e-22 wb0=8.421383269e-22 pb0=-1.612576997e-28 b1=4.817237160e-17 lb1=-9.224334748e-24 wb1=-4.145868451e-23 pb1=7.938757663e-30 keta=-3.217029525e-01 lketa=4.567993362e-08 wketa=2.835848705e-07 pketa=-5.430253251e-14 dwg=0.0 dwb=0.0 pclm=1.347544975e+00 lpclm=-2.123531822e-07 wpclm=-5.570907387e-07 ppclm=1.066750773e-13 pdiblc1=1.442850205e+00 lpdiblc1=-2.079304454e-07 wpdiblc1=-1.261081142e-06 ppdiblc1=2.414793836e-13 pdiblc2=1.734326396e-02 lpdiblc2=-1.711339459e-09 wpdiblc2=-1.802687858e-08 ppdiblc2=3.451894870e-15 pdiblcb=9.699306851e-01 lpdiblcb=-2.055078410e-07 wpdiblcb=-8.046569335e-07 ppdiblcb=1.540805376e-13 drout=1.380425306e+00 ldrout=-1.679521108e-07 wdrout=-1.154523721e-12 pdrout=2.206056431e-19 pscbe1=5.683221331e+09 lpscbe1=-9.367114926e+02 wpscbe1=-4.197000560e+03 ppscbe1=8.036668493e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.194670317e-05 lalpha0=9.951202500e-12 walpha0=4.473835125e-11 palpha0=-8.566767926e-18 alpha1=0.85 beta0=-4.234398384e+01 lbeta0=1.085035961e-05 wbeta0=4.806771689e-05 pbeta0=-9.204294837e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=3.936597724e+00 lkt1=-5.587614972e-07 wkt1=-3.640634028e-06 pkt1=4.895611021e-13 kt2=-3.712470563e-02 lkt2=1.578948873e-09 wkt2=-4.258501446e-09 pkt2=8.154434051e-16 at=5.967723227e+05 lat=-1.087739738e-01 wat=-4.563442222e-01 pat=8.738352974e-8 ute=-2.184033994e-02 lute=-2.483961869e-07 wute=-9.749215045e-07 pute=1.866838192e-13 ua1=5.468053699e-09 lua1=-1.051622161e-15 wua1=-3.028156686e-15 pua1=5.798496106e-22 ub1=-2.385362506e-18 lub1=5.922883493e-25 wub1=5.532839330e-25 pub1=-1.059461279e-31 uc1=4.059564858e-10 luc1=-4.955087738e-17 wuc1=-3.868236907e-16 puc1=7.407132126e-23 kt1l=0.0 prt=0.0 tvoff=1.654366268e-02 ltvoff=-2.275064842e-09 wtvoff=-1.258363923e-08 ptvoff=1.730487121e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.79 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='8.895100663e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-7.176191915e-09 wvth0=-2.254696290e-07 pvth0=-1.516550710e-14 k1=9.070734928e-01 lk1=-3.417968131e-16 wk1=-2.421362666e-15 pk1=2.941613619e-22 k2=-3.498052196e-01 lk2=4.798109350e-08 wk2=1.450533382e-07 pk2=-3.301736425e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587037853e-01 ldsub=-1.412889074e-11 wdsub=-5.612345314e-11 pdsub=1.074688124e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000028e-03 lcdscd=-3.616802170e-18 wcdscd=-2.429080548e-17 pcdscd=3.112735764e-24 cit=0.0 voff='-1.942012799e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.805764590e-08 wvoff=1.379748028e-06 pvoff=-8.192899335e-14 nfactor=-2.505169581e+01 lnfactor=2.168637153e-06 wnfactor=2.358661804e-05 pnfactor=-1.902404453e-12 eta0=-8.469097032e-03 leta0=1.754631528e-09 weta0=7.886176835e-09 peta0=-1.510092390e-15 etab=-4.399799988e-02 letab=-1.475794487e-17 wetab=-1.045483700e-16 petab=1.270115957e-23 u0=5.617407789e-02 lu0=-8.057028180e-09 wu0=-2.049849589e-08 pu0=6.184758901e-15 ua=-1.250950752e-09 lua=5.372357607e-17 wua=2.292405273e-17 pua=-3.525741114e-23 ub=2.937153980e-18 lub=-1.675648050e-25 wub=-6.253029444e-25 pub=1.471135007e-31 uc=-3.761214224e-10 luc=8.974593083e-17 wuc=3.770293721e-16 puc=-7.219584632e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.057378644e+05 lvsat=1.185258296e-03 wvsat=2.085862456e-02 pvsat=1.600100967e-10 a0=1.500000009e+00 la0=-1.044125675e-15 wa0=-7.396806723e-15 pa0=8.986082989e-22 ags=1.250000002e+00 lags=-2.235571728e-16 wags=-1.583721598e-15 pags=1.924003179e-22 a1=0.0 a2=0.42385546 b0=4.833567126e-07 lb0=-9.255604347e-14 wb0=-4.159922543e-13 pb0=7.965669280e-20 b1=-6.907728526e-10 lb1=1.322733305e-16 wb1=5.945012217e-16 pb1=-1.138386609e-22 keta=-1.356960822e-03 lketa=-1.566183894e-08 wketa=-1.363331660e-07 pketa=2.610589263e-14 dwg=0.0 dwb=0.0 pclm=1.084829369e+00 lpclm=-1.620468215e-07 wpclm=-5.656456552e-07 ppclm=1.083132240e-13 pdiblc1=3.569721485e-01 lpdiblc1=1.787521242e-16 wpdiblc1=1.266317717e-15 ppdiblc1=-1.538398298e-22 pdiblc2=8.406112139e-03 lpdiblc2=-4.792753000e-18 wpdiblc2=-3.395286829e-17 ppdiblc2=4.124797726e-24 pdiblcb=-1.032957699e-01 lpdiblcb=-1.419098172e-17 wpdiblcb=-1.005320271e-16 ppdiblcb=1.221323043e-23 drout=5.033266678e-01 ldrout=-9.467460149e-16 wdrout=-6.706946110e-15 pdrout=8.147997832e-22 pscbe1=7.914198808e+08 lpscbe1=-9.353065491e-08 wpscbe1=-6.625900269e-07 ppscbe1=8.049535751e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.324873625e-07 lalpha0=-2.123337781e-14 walpha0=-9.543321256e-14 palpha0=1.827412441e-20 alpha1=0.85 beta0=1.187370016e+01 lbeta0=4.684321719e-07 wbeta0=2.463837317e-06 pbeta0=-4.717903528e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=8.282568017e-01 lkt1=3.644227266e-08 wkt1=-9.202028314e-07 pkt1=-3.136338601e-14 kt2=-2.887893895e-02 lkt2=-5.673100878e-18 wkt2=-4.018951838e-17 pkt2=4.882455551e-24 at=-1.192221095e+05 lat=2.832893603e-02 wat=7.952768054e-02 pat=-1.522843743e-8 ute=-1.275698598e+00 lute=-8.299884468e-09 wute=-3.730375142e-08 pute=7.143146169e-15 ua1=-2.384732719e-11 lua1=-1.070419844e-24 wua1=-7.583076005e-24 pua1=9.212375687e-31 ub1=7.077531825e-19 lub1=-1.520583321e-33 wub1=-1.077212523e-32 pub1=1.308662271e-39 uc1=1.471862498e-10 luc1=2.201701467e-26 wuc1=1.559731763e-25 puc1=-1.894853648e-32 kt1l=0.0 prt=0.0 tvoff=9.220847822e-03 ltvoff=-8.728483167e-10 wtvoff=-7.013671921e-09 ptvoff=6.639163608e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.80 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='2.311839512e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.799693069e-07 wvth0=-1.383366554e-06 pvth0=1.255027587e-13 k1=0.90707349 k2=3.314829148e-01 lk2=-3.478587680e-08 wk2=-4.634451343e-07 pk2=4.090668119e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.584578332e-01 ldsub=1.575085221e-11 wdsub=1.309555803e-10 pdsub=-1.198060222e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999994e-03 lcdscd=5.364814495e-19 wcdscd=5.131929603e-18 pcdscd=-4.617131330e-25 cit=0.0 voff='-3.811502193e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.251744344e-07 wvoff=2.975917916e-06 pvoff=-2.758412884e-13 nfactor=-3.360042571e+01 lnfactor=3.207188154e-06 wnfactor=3.027358065e-05 pnfactor=-2.714776793e-12 eta0=2.419182927e-02 leta0=-2.213213472e-09 weta0=-1.840107703e-08 peta0=1.683440933e-15 etab=-0.043998 u0=-7.877763114e-02 lu0=8.337715144e-09 wu0=9.922485193e-08 pu0=-8.359951732e-15 ua=7.015588068e-10 lua=-1.834790002e-16 wua=-1.454022025e-15 pua=1.441708601e-22 ub=1.206464119e-18 lub=4.268978344e-26 wub=1.124571851e-24 pub=-6.547178873e-32 uc=1.233588525e-09 luc=-1.058112919e-16 wuc=-8.797352007e-16 puc=8.048345457e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.996883088e+04 lvsat=2.253116188e-02 wvsat=1.969530383e-01 pvsat=-2.123299586e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-8.616127790e-06 lb0=1.012903931e-12 wb0=5.917655792e-12 pb0=-6.897928737e-19 b1=1.231344836e-08 lb1=-1.447557488e-15 wb1=-8.457020513e-15 pb1=9.857945085e-22 keta=-4.452189562e-01 lketa=3.826117942e-08 wketa=3.181107210e-07 pketa=-2.910267742e-14 dwg=0.0 dwb=0.0 pclm=-8.461799054e-01 lpclm=7.254377113e-08 wpclm=8.439858005e-07 ppclm=-6.293726303e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.627532697e-07 lalpha0=2.678282563e-14 walpha0=2.226775051e-13 palpha0=-2.037187423e-20 alpha1=0.85 beta0=1.886497129e+01 lbeta0=-3.809093927e-07 wbeta0=-4.039363630e-06 pbeta0=3.182575176e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=5.404344724e+00 lkt1=-5.194883447e-07 wkt1=-4.858530532e-06 pkt1=4.470882931e-13 kt2=-0.028878939 at=2.976815455e+05 lat=-2.231902140e-02 wat=-1.855645879e-01 pat=1.697656189e-8 ute=-2.069266193e+00 lute=8.810746842e-08 wute=5.144396167e-07 pute=-5.988594865e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=8.680193499e-03 ltvoff=-8.071663855e-10 wtvoff=-7.999349171e-09 ptvoff=7.836623473e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.81 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.82 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.139140924e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.860518861e-06 wvth0=5.382371281e-08 pvth0=-1.073324816e-12 k1=7.676632329e-01 lk1=-3.981427614e-06 wk1=-1.042992115e-07 pk1=2.079881265e-12 k2=-1.386150690e-01 lk2=1.883956396e-06 wk2=5.176825013e-08 pk2=-1.032335835e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.900746404e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.235710083e-06 wvoff=4.571416589e-08 pvoff=-9.116083991e-13 nfactor=2.985057968e+00 lnfactor=-4.798878092e-06 wnfactor=-1.563755244e-07 pnfactor=3.118360330e-12 eta0=0.08 etab=-0.07 u0=1.990891099e-02 lu0=1.241973497e-07 wu0=3.062994800e-09 pu0=-6.108066793e-14 ua=-1.856302845e-09 lua=1.599803212e-14 wua=4.121610589e-16 pua=-8.219103986e-21 ub=2.761221281e-18 lub=-1.851150758e-23 wub=-5.424193951e-25 pub=1.081664877e-29 uc=6.614414220e-11 luc=-3.511125797e-16 wuc=-1.946723367e-18 puc=3.882055676e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.290558324e+00 la0=1.436618075e-06 wa0=6.722009529e-08 pa0=-1.340468589e-12 ags=5.067051857e-01 lags=-3.227034675e-06 wags=-1.245602882e-07 pags=2.483917243e-12 a1=0.0 a2=0.42385546 b0=4.881764970e-07 lb0=-8.296326155e-12 wb0=-2.801331174e-13 pb0=5.586270638e-18 b1=1.483684889e-07 lb1=-2.449183178e-12 wb1=-8.055833863e-14 pb1=1.606452982e-18 keta=-3.539403766e-02 lketa=6.151437463e-07 wketa=2.194674521e-08 pketa=-4.376507124e-13 dwg=0.0 dwb=0.0 pclm=-1.586863030e-01 lpclm=3.500953265e-06 wpclm=9.998431226e-08 ppclm=-1.993835763e-12 pdiblc1=0.39 pdiblc2=-8.256848595e-03 lpdiblc2=1.838041873e-07 wpdiblc2=5.908456205e-09 ppdiblc2=-1.178233967e-13 pdiblcb=1.224375199e+01 lpdiblcb=-2.446571460e-04 wpdiblcb=-8.227817682e-06 ppdiblcb=1.640749111e-10 drout=0.56 pscbe1=-5.566899859e+08 lpscbe1=1.558805991e+04 wpscbe1=3.245086203e+02 ppscbe1=-6.471184108e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.757351227e-01 lkt1=-2.122746707e-07 wkt1=-5.026222180e-09 pkt1=1.002303392e-13 kt2=-3.507328862e-02 lkt2=1.107820862e-07 wkt2=-2.450658404e-10 pkt2=4.886977025e-15 at=1.981626675e+05 lat=-4.618980097e-01 wat=-2.328306437e-16 ute=-8.899258942e-01 lute=-4.496288724e-06 wute=-8.477061289e-08 pute=1.690451990e-12 ua1=4.961274389e-10 lua1=1.246088743e-14 wua1=3.582121031e-16 pua1=-7.143281640e-21 ub1=1.285679393e-19 lub1=-1.391991379e-23 wub1=-3.433960004e-25 pub1=6.847826535e-30 uc1=9.616896630e-11 luc1=-1.243363703e-15 wuc1=-1.811577255e-17 puc1=3.612554246e-22 kt1l=0.0 prt=0.0 tvoff=9.855170968e-03 ltvoff=-1.447965451e-07 wtvoff=-5.478957267e-09 ptvoff=1.092585496e-13 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.83 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.452026980e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.374363673e-08 wvth0=-8.363868462e-08 pvth0=1.833088920e-14 k1=6.024347140e-01 lk1=-2.669267645e-06 wk1=-1.106043611e-07 pk1=2.129953523e-12 k2=-2.641305672e-02 lk2=9.929056862e-07 wk2=2.430771357e-08 pk2=-8.142583686e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.410326741e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.420532059e-07 wvoff=-1.442776698e-07 pvoff=5.972091045e-13 nfactor=5.752657252e-01 lnfactor=1.433845327e-05 wnfactor=1.573601050e-06 pnfactor=-1.062022441e-11 eta0=0.08 etab=-0.07 u0=5.246237643e-02 lu0=-1.343255403e-07 wu0=-1.688778591e-08 pu0=9.735817777e-14 ua=1.991936389e-09 lua=-1.456270589e-14 wua=-1.990084035e-15 pua=1.085829179e-20 ub=-9.537389584e-19 lub=1.099079715e-23 wub=1.872737418e-24 pub=-8.363285241e-30 uc=1.489389182e-10 luc=-1.008626134e-15 wuc=-9.334787111e-17 puc=7.646814920e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.944146108e+00 la0=-3.753840160e-06 wa0=-3.590984031e-07 pa0=2.045133798e-12 ags=2.239821887e-01 lags=-9.817939522e-07 wags=9.198571050e-08 pags=7.642202259e-13 a1=0.0 a2=0.42385546 b0=-2.897096051e-07 lb0=-2.118754566e-12 wb0=2.203623963e-13 pb0=1.611592523e-18 b1=-1.004745941e-09 lb1=-1.262937724e-12 wb1=7.642419143e-16 pb1=9.606308471e-19 keta=2.246824877e-02 lketa=1.556312086e-07 wketa=-2.672087318e-08 pketa=-5.115750228e-14 dwg=0.0 dwb=0.0 pclm=2.088219555e+00 lpclm=-1.434281815e-05 wpclm=-1.861829491e-06 ppclm=1.358588109e-11 pdiblc1=0.39 pdiblc2=3.704385420e-02 lpdiblc2=-1.759507098e-07 wpdiblc2=-2.592607222e-08 ppdiblc2=1.349900651e-13 pdiblcb=-3.683125596e+01 lpdiblcb=1.450713426e-04 wpdiblcb=2.468345305e-05 ppdiblcb=-9.728948462e-11 drout=0.56 pscbe1=1.807620282e+09 lpscbe1=-3.188076984e+03 wpscbe1=-7.834961505e+02 ppscbe1=2.328020267e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.281997972e-01 lkt1=2.043728068e-07 wkt1=2.809151204e-08 pkt1=-1.627736834e-13 kt2=-1.002079484e-01 lkt2=6.280480747e-07 wkt2=6.057073523e-08 pkt2=-4.780808558e-13 at=140000.0 ute=-3.391837737e+00 lute=1.537260915e-05 wute=1.448924565e-06 pute=-1.048936679e-11 ua1=-6.876590069e-10 lua1=2.186191092e-14 wua1=1.476272352e-15 pua1=-1.602234145e-20 ub1=-2.654941034e-19 lub1=-1.079047560e-23 wub1=-5.099632445e-25 pub1=8.170617972e-30 uc1=2.699318853e-10 luc1=-2.623299491e-15 wuc1=-2.284741847e-16 puc1=2.031813810e-21 kt1l=0.0 prt=0.0 tvoff=-1.701995802e-02 ltvoff=6.863191557e-08 wtvoff=1.530425160e-08 ptvoff=-5.579101263e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.84 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.225817059e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.129039605e-07 wvth0=-6.240820053e-08 pvth0=-6.534876661e-14 k1=-4.274317175e-01 lk1=1.389936476e-06 wk1=6.617152121e-07 pk1=-9.141332624e-13 k2=3.071412381e-01 lk2=-3.217938970e-07 wk2=-2.298068179e-07 pk2=1.873304997e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.610037732e+00 ldsub=8.553173340e-06 wdsub=1.650600140e-06 pdsub=-6.505817344e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.809953163e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.903924111e-07 wvoff=-4.537024033e-08 pvoff=2.073668557e-13 nfactor=6.438542122e+00 lnfactor=-8.771568564e-06 wnfactor=-2.745144208e-06 pnfactor=6.402049557e-12 eta0=-4.950599990e-01 leta0=2.266590935e-06 weta0=4.374090371e-07 peta0=-1.724041596e-12 etab=4.327254079e-01 letab=-1.981485157e-06 wetab=-3.823890325e-07 petab=1.507181018e-12 u0=3.087130085e-02 lu0=-4.922461815e-08 wu0=-7.424603310e-10 pu0=3.372160304e-14 ua=3.086947559e-09 lua=-1.887867708e-14 wua=-2.540049415e-15 pua=1.302597264e-20 ub=-5.055025882e-18 lub=2.715596214e-23 wub=4.565269925e-24 pub=-1.897586442e-29 uc=-2.872034573e-10 luc=7.104229331e-16 wuc=2.165546920e-16 puc=-4.567951218e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=-9.484906727e-01 la0=7.647447213e-06 wa0=1.711735117e-06 pa0=-6.117027531e-12 ags=-3.383542104e-01 lags=1.234647092e-06 wags=4.469404682e-07 pags=-6.348289820e-13 a1=0.0 a2=0.42385546 b0=-6.740571655e-07 lb0=-6.038540378e-13 wb0=5.127094499e-13 pb0=4.593107045e-19 b1=-3.861297578e-07 lb1=2.550271184e-13 wb1=2.937026500e-13 pb1=-1.939817871e-19 keta=2.309594397e-01 lketa=-6.661339017e-07 wketa=-1.545151428e-07 pketa=4.525418222e-13 dwg=0.0 dwb=0.0 pclm=-3.969017693e+00 lpclm=9.531697662e-06 wpclm=3.406831033e-06 ppclm=-7.180470602e-12 pdiblc1=0.39 pdiblc2=-6.491634393e-03 lpdiblc2=-4.356190977e-09 wpdiblc2=6.040269373e-09 ppdiblc2=8.995177269e-15 pdiblcb=6.541823883e-02 lpdiblcb=-3.563822225e-07 wpdiblcb=-6.877500584e-08 ppdiblcb=2.710757227e-13 drout=0.56 pscbe1=1.191722126e+09 lpscbe1=-7.605230234e+02 wpscbe1=-3.800594207e+02 ppscbe1=7.378800444e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-5.662826980e-01 lkt1=1.142773227e-06 wkt1=2.058286087e-07 pkt1=-8.633219615e-13 kt2=-8.737585318e-02 lkt2=5.774705511e-07 wkt2=4.850218503e-08 pkt2=-4.305128341e-13 at=1.547201682e+05 lat=-5.801933702e-02 wat=1.006866085e-02 pat=-3.968548580e-8 ute=-8.048884277e+00 lute=3.372829289e-05 wute=4.807006019e-06 pute=-2.372519783e-11 ua1=-2.118006063e-08 lua1=1.026324250e-13 wua1=1.562597908e-14 pua1=-7.179321241e-20 ub1=1.762162534e-17 lub1=-8.129230647e-23 wub1=-1.280468812e-23 pub1=5.663010393e-29 uc1=-1.224678124e-10 luc1=-1.076661576e-15 wuc1=8.805719376e-17 puc1=7.842098130e-22 kt1l=0.0 prt=0.0 tvoff=-1.576789054e-03 ltvoff=7.762881285e-09 wtvoff=3.264733805e-09 ptvoff=-8.337421787e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.85 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.547453489e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.446072979e-07 wvth0=-1.406525128e-08 pvth0=-1.592059258e-13 k1=6.344675071e-01 lk1=-6.717260016e-07 wk1=-2.921618237e-08 pk1=4.273003670e-13 k2=9.579544350e-02 lk2=8.853100431e-08 wk2=-1.137933118e-07 pk2=-3.790809831e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.182521264e+00 ldsub=-4.634484855e-06 wdsub=-3.301200280e-06 pdsub=3.108033847e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.124977389e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.292308986e-07 wvoff=2.337032585e-08 pvoff=7.390800887e-14 nfactor=2.364783560e+00 lnfactor=-8.624233484e-07 wnfactor=5.371591555e-07 pnfactor=2.950352930e-14 eta0=1.303055344e+00 leta0=-1.224424829e-06 weta0=-8.748178074e-07 peta0=8.236284515e-13 etab=-1.061916955e+00 letab=9.203420646e-07 wetab=7.647780649e-07 petab=-7.200278412e-13 u0=8.739506644e-04 lu0=9.014817263e-09 wu0=2.159806098e-08 pu0=-9.652206314e-15 ua=-9.794342704e-09 lua=6.130167626e-15 wua=6.737725380e-15 pua=-4.986697234e-21 ub=1.399120584e-17 lub=-9.822030090e-24 wub=-9.141592746e-24 pub=7.635817555e-30 uc=-1.278278308e-10 luc=4.009973853e-16 wuc=1.268817697e-16 puc=-2.826963986e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.439540702e+04 lvsat=1.079555388e-01 wvsat=3.513338898e-02 pvsat=-6.821098283e-8 a0=7.714141406e+00 la0=-9.170931691e-06 wa0=-4.831070121e-06 pa0=6.585737240e-12 ags=4.826954050e+00 lags=-8.793726582e-06 wags=-3.405999461e-06 pags=6.845599950e-12 a1=0.0 a2=0.42385546 b0=-1.538230396e-07 lb0=-1.613881310e-12 wb0=1.170027263e-13 pb0=1.227569768e-18 b1=-3.849097230e-07 lb1=2.526584378e-13 wb1=2.927746524e-13 pb1=-1.921800929e-19 keta=-7.333499124e-01 lketa=1.206059205e-06 wketa=5.379187702e-07 pketa=-8.918089258e-13 dwg=0.0 dwb=0.0 pclm=2.454893794e+00 lpclm=-2.940236555e-06 wpclm=-1.537500137e-06 ppclm=2.418879142e-12 pdiblc1=5.481820911e-01 lpdiblc1=-3.071083154e-07 wpdiblc1=-8.358448819e-08 ppdiblc1=1.622781136e-13 pdiblc2=-3.022798571e-02 lpdiblc2=4.172760279e-08 wpdiblc2=2.665632377e-08 ppdiblc2=-3.103060371e-14 pdiblcb=1.621371179e-01 lpdiblcb=-5.441605722e-07 wpdiblcb=-1.248887102e-07 ppdiblcb=3.800196941e-13 drout=4.378077866e+00 ldrout=-7.412744724e-06 wdrout=-2.787638631e-06 pdrout=5.412161375e-12 pscbe1=3.362586588e+08 lpscbe1=9.003473216e+02 wpscbe1=3.527365039e+02 ppscbe1=-6.848329839e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.855437731e-05 lalpha0=-7.479453921e-11 walpha0=-2.930201482e-11 palpha0=5.688945154e-17 alpha1=2.067411445e+00 lalpha1=-2.363587276e-06 walpha1=-8.164350719e-07 palpha1=1.585097262e-12 beta0=3.914368737e+01 lbeta0=-4.908792506e-05 wbeta0=-1.923158169e-05 pbeta0=3.733784662e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=1.585687332e-01 lkt1=-2.645156786e-07 wkt1=-3.675665927e-07 pkt1=2.499167944e-13 kt2=5.057860012e-01 lkt2=-5.741448849e-07 wkt2=-3.849108965e-07 pkt2=4.109525959e-13 at=1.236387502e+02 lat=2.421276606e-01 wat=1.027386646e-01 pat=-2.196030007e-7 ute=1.889194669e+01 lute=-1.857695326e-05 wute=-1.424406546e-05 pute=1.326219074e-11 ua1=6.058564990e-08 lua1=-5.611455725e-14 wua1=-4.164376561e-14 pua1=3.939519512e-20 ub1=-4.567435484e-17 lub1=4.159595291e-23 wub1=3.125045807e-23 pub1=-2.890234563e-29 uc1=-1.170285928e-09 luc1=9.576626256e-16 wuc1=8.326064145e-16 puc1=-6.613220754e-22 kt1l=0.0 prt=0.0 tvoff=3.794700004e-03 ltvoff=-2.665789521e-09 wtvoff=-1.957738162e-09 ptvoff=1.801934423e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.86 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.086730622e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.562493888e-07 wvth0=-3.448963259e-07 pvth0=1.522668993e-13 k1=-5.681650689e-01 lk1=4.605357319e-07 wk1=7.995874806e-07 pk1=-3.530066785e-13 k2=3.693794794e-01 lk2=-1.690445353e-07 wk2=-2.900858165e-07 pk2=1.280688268e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-7.200593438e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.544826465e-07 wvoff=1.918216869e-07 pvoff=-8.468658928e-14 nfactor=-1.608530620e+00 lnfactor=2.878396325e-06 wnfactor=1.070462708e-06 pnfactor=-4.725942991e-13 eta0=-4.278892114e-01 leta0=4.052352364e-07 weta0=-5.336176943e-13 peta0=2.355847411e-19 etab=-1.583239050e-01 letab=6.962185878e-8 u0=-1.902015903e-03 lu0=1.162835092e-08 wu0=2.136413145e-08 pu0=-9.431964935e-15 ua=-4.902847280e-09 lua=1.524893165e-15 wua=2.713553765e-15 pua=-1.197995997e-21 ub=4.804488238e-18 lub=-1.172864086e-24 wub=-1.941728065e-24 pub=8.572457565e-31 uc=5.149098445e-10 luc=-2.041311376e-16 wuc=-3.264779776e-16 puc=1.441354564e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.408780160e+05 lvsat=-1.711206813e-03 wvsat=-7.026677795e-02 pvsat=3.102179873e-8 a0=-5.038914142e+00 la0=2.835891564e-06 wa0=4.074704712e-06 pa0=-1.798925084e-12 ags=-8.636398218e+00 lags=3.881831091e-06 wags=7.277798282e-06 pags=-3.213046052e-12 a1=0.0 a2=0.42385546 b0=-3.517407096e-06 lb0=1.552885989e-12 wb0=2.675452394e-12 pb0=-1.181174776e-18 b1=-2.194573553e-07 lb1=9.688734994e-14 wb1=1.669262871e-13 pb1=-7.369561876e-20 keta=1.037521915e+00 lketa=-4.611918285e-07 wketa=-7.707318690e-07 pketa=3.402673299e-13 dwg=0.0 dwb=0.0 pclm=-1.656912412e+00 lpclm=9.309714225e-07 wpclm=1.942688577e-06 ppclm=-8.576698091e-13 pdiblc1=3.888287494e-01 lpdiblc1=-1.570793751e-07 wpdiblc1=1.671689764e-07 ppdiblc1=-7.380276271e-14 pdiblc2=2.649575172e-02 lpdiblc2=-1.167700187e-08 wpdiblc2=-1.186809615e-08 ppdiblc2=5.239598297e-15 pdiblcb=-6.994877397e-01 lpdiblcb=2.670471685e-07 wpdiblcb=5.248774438e-07 ppdiblcb=-2.317260432e-13 drout=-7.464663324e+00 ldrout=3.737030308e-06 wdrout=5.575277262e-06 pdrout=-2.461406857e-12 pscbe1=2.048048307e+09 lpscbe1=-7.112786670e+02 wpscbe1=-7.054730077e+02 ppscbe1=3.114564563e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.043585627e-05 lalpha0=3.723309984e-11 walpha0=5.860402963e-11 palpha0=-2.587285863e-17 alpha1=-1.584822889e+00 lalpha1=1.074940218e-06 walpha1=1.632870144e-06 palpha1=-7.208893083e-13 beta0=-4.037877232e+01 lbeta0=2.578135742e-05 wbeta0=3.846316339e-05 pbeta0=-1.698094815e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=3.501116764e-01 lkt1=-4.448506780e-07 wkt1=-1.922840133e-07 pkt1=8.489069990e-14 kt2=-1.634873959e-01 lkt2=5.596664860e-08 wkt2=9.712875115e-08 pkt2=-4.288098383e-14 at=4.750798333e+05 lat=-2.050369471e-01 wat=-2.457519726e-01 pat=1.084960554e-7 ute=-4.239603029e-01 lute=-3.912972522e-07 wute=-2.967949597e-07 pute=1.310308196e-13 ua1=1.117626906e-09 lua1=-1.262461602e-16 wua1=3.763456183e-16 pua1=-1.661513216e-22 ub1=-2.253694004e-18 lub1=7.160086188e-25 wub1=1.039046286e-24 pub1=-4.587243888e-31 uc1=-2.933590204e-10 luc1=1.320482191e-16 wuc1=2.451304148e-16 puc1=-1.082216463e-22 kt1l=0.0 prt=0.0 tvoff=1.813734813e-03 ltvoff=-8.007385278e-10 wtvoff=-8.249729550e-11 ptvoff=3.642140100e-17 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.87 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.482941075e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.853720580e-8 k1=1.440277360e-01 lk1=1.461125792e-7 k2=7.969704024e-02 lk2=-4.115379395e-08 pk2=1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-1.169482067e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.178247696e-8 nfactor=5.439654304e+00 lnfactor=-2.332786435e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 wetab=1.214306433e-23 petab=4.336808690e-31 u0=2.047379937e-02 lu0=1.749741742e-9 ua=-1.652990168e-09 lua=9.012674784e-17 ub=2.069596195e-18 lub=3.455246251e-26 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.343617910e+05 lvsat=1.165615310e-3 a0=1.296210063e+00 la0=3.902291978e-8 ags=-6.815012482e-01 lags=3.698554480e-07 pags=-1.665334537e-28 a1=0.0 a2=0.42385546 b0=1.286445378e-16 lb0=-2.463362796e-23 b1=-6.333203389e-18 lb1=1.212719784e-24 keta=5.112499917e-02 lketa=-2.571139952e-08 wketa=1.387778781e-23 pketa=-1.734723476e-30 dwg=0.0 dwb=0.0 pclm=6.151398981e-01 lpclm=-7.210786349e-8 pdiblc1=-2.150883798e-01 lpdiblc1=1.095415826e-07 wpdiblc1=5.551115123e-23 ppdiblc1=4.163336342e-29 pdiblc2=-6.356604809e-03 lpdiblc2=2.826853610e-09 wpdiblc2=-4.336808690e-25 ppdiblc2=-5.014435048e-31 pdiblcb=-8.794872769e-02 lpdiblcb=-2.938743745e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406427e+08 lpscbe1=1.198662602e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637210e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-8.497299977e-01 lkt1=8.486262334e-8 kt2=-4.272334130e-02 lkt2=2.651009219e-9 at=-3.181692162e+03 lat=6.108820679e-03 pat=-3.637978807e-24 ute=-1.303565937e+00 lute=-2.963679149e-9 ua1=1.486947612e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 pub1=1.925929944e-46 uc1=-1.025991505e-10 luc1=4.783040721e-17 wuc1=-4.523643975e-32 puc1=-1.615587134e-39 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.88 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493605488e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810552122e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.754989805e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940211880e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372706393e-16 ags=1.250000000e+00 lags=2.939115618e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-8 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350031281e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301036082e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865674282e-18 drout=5.033266590e-01 ldrout=1.244684356e-16 pscbe1=7.914198799e+08 lpscbe1=1.229619980e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458339502e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407276948e-25 ub1=7.077531684e-19 lub1=1.999107579e-34 uc1=1.471862500e-10 luc1=-2.894511758e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.89 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-9.079060523e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.552352942e-07 wvth0=1.065674954e-06 pvth0=-1.294645874e-13 k1=0.90707349 k2=-9.580463684e-01 lk2=1.016335849e-07 wk2=5.174121035e-07 pk2=-6.285832680e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999998e-03 lcdscd=2.111323269e-19 wcdscd=1.763506008e-18 pcdscd=-2.142418187e-25 cit=0.0 voff='2.399373771e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.167023115e-07 wvoff=-1.748273090e-06 pvoff=2.123907046e-13 nfactor=1.471786983e+01 lnfactor=-1.396704025e-06 wnfactor=-6.478861125e-06 pnfactor=7.870909227e-13 eta0=8.115409484e-10 leta0=-7.424687366e-17 weta0=-5.702435093e-20 peta0=6.927660297e-27 etab=-0.043998 u0=2.183619187e-01 lu0=-2.290346319e-08 wu0=-1.267889981e-07 pu0=1.540308823e-14 ua=-1.581850071e-09 lua=5.123179138e-17 wua=2.828118361e-16 pua=-3.435767872e-23 ub=5.346041977e-18 lub=-3.666730364e-25 wub=-2.024123534e-24 pub=2.459026716e-31 uc=7.700399989e-11 luc=9.689386900e-27 wuc=-1.209751646e-28 puc=1.470830527e-35 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.506710915e+05 lvsat=-2.502885432e-02 wvsat=-1.229991471e-01 pvsat=1.494267438e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-7.340024972e-06 lb0=8.961585444e-13 wb0=4.947011153e-12 pb0=-6.009925969e-19 b1=1.048972263e-08 lb1=-1.280711538e-15 wb1=-7.069836362e-15 pb1=8.588861403e-22 keta=-2.700000006e-02 lketa=5.207917431e-18 wketa=6.905587213e-20 pketa=-8.403000518e-27 dwg=0.0 dwb=0.0 pclm=8.890083817e-01 lpclm=-8.620165949e-08 wpclm=-4.758539367e-07 ppclm=5.780959135e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.163942384e-24 walpha0=-1.382781286e-25 palpha0=1.680831005e-32 alpha1=0.85 beta0=1.125417800e+01 lbeta0=3.169516113e-07 wbeta0=1.749649290e-06 pbeta0=-2.125578936e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-4.852034439e+00 lkt1=5.383126064e-07 wkt1=2.942799664e-06 pkt1=-3.575089600e-13 kt2=-0.028878939 at=5.372048694e+04 lat=5.715526640e-12 wat=-2.933666110e-14 pat=3.579771146e-21 ute=-1.967998703e+00 lute=7.923790317e-08 wute=4.374123232e-07 pute=-5.313947349e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-1.552129144e-02 ltvoff=1.885619612e-09 wtvoff=1.040907472e-08 ptvoff=-1.264556852e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.90 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.91 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-7 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-08 wu0=-2.220446049e-22 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 uc=6.324132312e-11 luc=-2.932260536e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 b1=2.824547271e-08 lb1=-5.375173124e-14 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-7 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-7 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.92 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-07 pk2=-8.881784197e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-7 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 uc=9.745036742e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-8 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=1.776356839e-21 ppclm=2.486899575e-26 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116797e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 wua1=1.323488980e-29 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 wuc1=-2.067951531e-31 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.93 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 wua=6.617444900e-30 ub=1.752388505e-18 lub=-1.139532890e-24 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929614e-08 lb1=-3.422509015e-14 wb1=4.235164736e-28 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-6 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-8 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-1 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 wua1=1.323488980e-29 pua1=-2.646977960e-35 ub1=-1.471838908e-18 lub1=3.150583117e-24 wub1=1.232595164e-38 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.94 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-8 k2=-7.388526331e-02 lk2=3.200507309e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-7 eta0=-1.412393437e-03 leta0=3.712885085e-09 weta0=-6.938893904e-24 peta0=-1.387778781e-29 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=-7.632783294e-23 petab=-2.914335440e-28 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-6 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=-1.110223025e-22 pketa=-4.440892099e-28 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-9 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=4.658681210e-27 palpha0=7.199780052e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-8 at=1.533204212e+05 lat=-8.532912747e-2 ute=-2.347817386e+00 lute=1.198707212e-6 ua1=-1.510649725e-09 lua1=2.628829754e-15 wua1=-6.617444900e-30 pua1=-1.654361225e-36 ub1=9.241642797e-19 lub1=-1.501223529e-24 wub1=1.540743956e-39 pub1=6.162975822e-45 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.95 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.724451032e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.919953230e-8 k1=6.241244142e-01 lk1=-6.584338284e-8 k2=-6.317640297e-02 lk2=2.192283100e-08 wk2=4.440892099e-22 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.340281270e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.282038687e-07 wvoff=-3.552713679e-21 nfactor=-1.233075445e-02 lnfactor=2.173696432e-6 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=4.718447855e-22 peta0=1.804112415e-28 etab=-1.583239050e-01 letab=6.962185878e-8 u0=2.995469753e-02 lu0=-2.435942066e-9 ua=-8.565838072e-10 lua=-2.614755107e-16 ub=1.909117804e-18 lub=1.054014256e-25 uc=2.808849156e-11 luc=1.079367420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.610106241e+04 lvsat=4.454635133e-2 a0=1.037003369e+00 la0=1.534590465e-7 ags=2.215750624e+00 lags=-9.092406921e-7 a1=0.0 a2=0.42385546 b0=4.720422506e-07 lb0=-2.084000450e-13 b1=2.945156506e-08 lb1=-1.300245365e-14 keta=-1.117400778e-01 lketa=4.619125186e-8 dwg=0.0 dwb=0.0 pclm=1.239890271e+00 lpclm=-3.479264068e-7 pdiblc1=6.380995512e-01 lpdiblc1=-2.671289443e-07 wpdiblc1=3.552713679e-21 pdiblc2=8.798868558e-03 lpdiblc2=-3.864075705e-9 pdiblcb=8.317315893e-02 lpdiblcb=-7.848666098e-08 wpdiblcb=-6.591949209e-23 ppdiblcb=6.071532166e-29 drout=8.488040648e-01 ldrout=6.675084449e-8 pscbe1=9.960958087e+08 lpscbe1=-2.468563664e+02 wpscbe1=7.629394531e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414640e-06 lalpha0=-1.346715357e-12 alpha1=0.85 beta0=1.697483351e+01 lbeta0=4.605433985e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=6.339107061e-02 lkt1=-3.182675446e-7 kt2=-1.865572788e-02 lkt2=-7.974505161e-9 at=1.086315090e+05 lat=-4.325514223e-2 ute=-8.665203951e-01 lute=-1.959131673e-7 ua1=1.678807431e-09 lua1=-3.739995058e-16 wua1=-1.323488980e-29 ub1=-7.043401311e-19 lub1=3.199057494e-26 uc1=7.216247987e-11 luc1=-2.932440595e-17 kt1l=0.0 prt=0.0 tvoff=1.690720559e-03 ltvoff=-7.464294566e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.96 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.482941075e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.853720580e-8 k1=1.440277360e-01 lk1=1.461125792e-7 k2=7.969704024e-02 lk2=-4.115379395e-08 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-1.169482067e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.178247696e-8 nfactor=5.439654304e+00 lnfactor=-2.332786435e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 wetab=-4.857225733e-23 petab=2.081668171e-29 u0=2.047379937e-02 lu0=1.749741742e-9 ua=-1.652990168e-09 lua=9.012674784e-17 ub=2.069596195e-18 lub=3.455246251e-26 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.343617910e+05 lvsat=1.165615310e-3 a0=1.296210063e+00 la0=3.902291978e-8 ags=-6.815012482e-01 lags=3.698554480e-07 pags=1.776356839e-27 a1=0.0 a2=0.42385546 b0=1.286445378e-16 lb0=-2.463362796e-23 b1=-6.333203389e-18 lb1=1.212719784e-24 keta=5.112499917e-02 lketa=-2.571139952e-08 wketa=-2.220446049e-22 pketa=-2.775557562e-29 dwg=0.0 dwb=0.0 pclm=6.151398981e-01 lpclm=-7.210786349e-8 pdiblc1=-2.150883798e-01 lpdiblc1=1.095415826e-07 ppdiblc1=-2.775557562e-28 pdiblc2=-6.356604809e-03 lpdiblc2=2.826853610e-09 wpdiblc2=-1.951563910e-23 ppdiblc2=5.963111949e-30 pdiblcb=-8.794872769e-02 lpdiblcb=-2.938743745e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406427e+08 lpscbe1=1.198662602e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637210e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-8.497299977e-01 lkt1=8.486262334e-8 kt2=-4.272334130e-02 lkt2=2.651009219e-9 at=-3.181692162e+03 lat=6.108820679e-3 ute=-1.303565937e+00 lute=-2.963679149e-9 ua1=1.486947612e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 wub1=-6.162975822e-39 uc1=-1.025991505e-10 luc1=4.783040721e-17 wuc1=-2.067951531e-31 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.97 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493116990e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810552122e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.755015826e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940225758e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372697511e-16 ags=1.250000000e+00 lags=2.939160026e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-08 wketa=-1.776356839e-21 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.349942463e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301070776e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865618771e-18 drout=5.033266590e-01 ldrout=1.244675474e-16 pscbe1=7.914198799e+08 lpscbe1=1.229858398e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458478279e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407277206e-25 ub1=7.077531684e-19 lub1=1.999115282e-34 uc1=1.471862500e-10 luc1=-2.894304963e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.98 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.263974810e+01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.490615018e-06 wvth0=-8.019815444e-06 pvth0=9.742952990e-13 k1=0.90707349 k2=5.190481676e+00 lk2=-6.453264930e-07 wk2=-3.605987556e-06 pk2=4.380770042e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000019e-03 lcdscd=-2.287316170e-18 wcdscd=-1.202854483e-17 pcdscd=1.461303301e-24 cit=0.0 voff='-2.215680733e+01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.666529906e-06 wvoff=1.471988775e-05 pvoff=-1.788260284e-12 nfactor=-4.643032663e+01 lnfactor=6.031945771e-06 wnfactor=3.452907617e-05 pnfactor=-4.194799347e-12 eta0=8.107679152e-10 leta0=-7.415295110e-17 weta0=4.614508521e-19 peta0=-5.605981822e-26 etab=-0.043998 u0=-1.133993735e+00 lu0=1.413888157e-07 wu0=7.801439785e-07 pu0=-9.477657137e-14 ua=7.021761111e-09 lua=-9.939865167e-16 wua=-5.487045138e-15 pua=6.665991657e-22 ub=-4.870249054e-18 lub=8.744632958e-25 wub=4.827248153e-24 pub=-5.864430691e-31 uc=7.700399989e-11 luc=9.860406492e-27 wuc=8.238718901e-28 puc=-1.000888541e-34 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-2.675112995e+06 lvsat=3.425615512e-01 wvsat=1.906188486e+00 pvsat=-2.315752144e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-7.340013816e-06 lb0=8.961571891e-13 wb0=4.947003672e-12 pb0=-6.009916881e-19 b1=1.048973181e-08 lb1=-1.280712653e-15 wb1=-7.069842518e-15 pb1=8.588868882e-22 keta=-2.700000006e-02 lketa=5.109801471e-18 wketa=-4.733990977e-19 pketa=5.745404152e-26 dwg=0.0 dwb=0.0 pclm=8.890083656e-01 lpclm=-8.620165753e-08 wpclm=-4.758539259e-07 ppclm=5.780959004e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-9.675233840e-25 walpha0=9.461358021e-25 palpha0=-1.148788435e-31 alpha1=0.85 beta0=1.121716203e+01 lbeta0=3.214485331e-07 wbeta0=1.774473382e-06 pbeta0=-2.155736733e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=3.497658117e+01 lkt1=-4.300306590e-06 wkt1=-2.376754448e-05 pkt1=2.887423909e-12 kt2=-0.028878939 at=5.372048694e+04 lat=5.757668987e-12 wat=2.011656761e-13 pat=-2.468004823e-20 ute=-1.977252686e+00 lute=8.036213247e-08 wute=4.436183399e-07 pute=-5.389341764e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=1.440432657e-01 ltvoff=-1.749924018e-08 wtvoff=-9.660002336e-08 ptvoff=1.173555044e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.99 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.100 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-07 wvoff=8.881784197e-22 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-8 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 uc=6.324132312e-11 luc=-2.932260536e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 wb0=-2.117582368e-28 b1=2.824547271e-08 lb1=-5.375173124e-14 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-07 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+03 ppscbe1=7.629394531e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-7 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 wuc1=-1.033975766e-31 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.101 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-07 pk2=-2.220446049e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-7 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 uc=9.745036741e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-08 pketa=-1.110223025e-28 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=4.440892099e-22 ppclm=7.105427358e-27 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116796e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-08 wtvoff=-1.387778781e-23 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.102 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 ub=1.752388505e-18 lub=-1.139532890e-24 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929613e-08 lb1=-3.422509015e-14 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-6 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-8 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-01 wat=4.656612873e-16 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 wua1=3.308722450e-30 ub1=-1.471838908e-18 lub1=3.150583117e-24 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-09 wtvoff=-6.938893904e-24 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.103 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-08 wk1=-1.776356839e-21 k2=-7.388526331e-02 lk2=3.200507309e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-7 eta0=-1.412393438e-03 leta0=3.712885085e-09 weta0=1.734723476e-24 peta0=1.734723476e-30 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=-3.642919300e-23 petab=8.153200337e-29 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 pua=1.654361225e-36 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-06 pags=-1.776356839e-27 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=2.775557562e-23 pketa=1.110223025e-28 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-9 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=-3.176373552e-27 palpha0=-5.188076802e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-8 at=1.533204212e+05 lat=-8.532912747e-2 ute=-2.347817386e+00 lute=1.198707212e-6 ua1=-1.510649725e-09 lua1=2.628829754e-15 wua1=-8.271806126e-31 pua1=-3.308722450e-36 ub1=9.241642797e-19 lub1=-1.501223529e-24 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.104 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.724451032e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.919953230e-8 k1=6.241244142e-01 lk1=-6.584338284e-8 k2=-6.317640297e-02 lk2=2.192283100e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.340281270e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.282038687e-7 nfactor=-1.233075445e-02 lnfactor=2.173696432e-6 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=3.608224830e-22 peta0=1.908195824e-28 etab=-1.583239050e-01 letab=6.962185878e-08 wetab=-4.440892099e-22 u0=2.995469753e-02 lu0=-2.435942066e-9 ua=-8.565838072e-10 lua=-2.614755107e-16 ub=1.909117804e-18 lub=1.054014256e-25 uc=2.808849156e-11 luc=1.079367420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.610106241e+04 lvsat=4.454635133e-2 a0=1.037003369e+00 la0=1.534590465e-7 ags=2.215750624e+00 lags=-9.092406921e-7 a1=0.0 a2=0.42385546 b0=4.720422506e-07 lb0=-2.084000450e-13 b1=2.945156506e-08 lb1=-1.300245365e-14 keta=-1.117400778e-01 lketa=4.619125186e-8 dwg=0.0 dwb=0.0 pclm=1.239890271e+00 lpclm=-3.479264068e-7 pdiblc1=6.380995512e-01 lpdiblc1=-2.671289443e-7 pdiblc2=8.798868558e-03 lpdiblc2=-3.864075705e-9 pdiblcb=8.317315893e-02 lpdiblcb=-7.848666098e-08 wpdiblcb=-1.214306433e-23 ppdiblcb=-2.255140519e-29 drout=8.488040648e-01 ldrout=6.675084449e-8 pscbe1=9.960958087e+08 lpscbe1=-2.468563664e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414640e-06 lalpha0=-1.346715357e-12 alpha1=0.85 beta0=1.697483351e+01 lbeta0=4.605433985e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=6.339107061e-02 lkt1=-3.182675446e-7 kt2=-1.865572788e-02 lkt2=-7.974505161e-9 at=1.086315090e+05 lat=-4.325514223e-2 ute=-8.665203951e-01 lute=-1.959131673e-7 ua1=1.678807431e-09 lua1=-3.739995058e-16 ub1=-7.043401311e-19 lub1=3.199057494e-26 uc1=7.216247987e-11 luc1=-2.932440595e-17 wuc1=2.067951531e-31 kt1l=0.0 prt=0.0 tvoff=1.690720559e-03 ltvoff=-7.464294566e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.105 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.482941075e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.853720580e-8 k1=1.440277360e-01 lk1=1.461125792e-7 k2=7.969704024e-02 lk2=-4.115379395e-08 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-1.169482067e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.178247696e-8 nfactor=5.439654304e+00 lnfactor=-2.332786435e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 wetab=1.734723476e-24 petab=1.084202172e-29 u0=2.047379937e-02 lu0=1.749741742e-9 ua=-1.652990168e-09 lua=9.012674784e-17 ub=2.069596195e-18 lub=3.455246251e-26 wub=6.162975822e-39 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.343617910e+05 lvsat=1.165615310e-3 a0=1.296210063e+00 la0=3.902291978e-8 ags=-6.815012482e-01 lags=3.698554480e-07 wags=-8.881784197e-22 pags=-1.110223025e-28 a1=0.0 a2=0.42385546 b0=1.286445378e-16 lb0=-2.463362796e-23 b1=-6.333203389e-18 lb1=1.212719784e-24 keta=5.112499917e-02 lketa=-2.571139952e-08 wketa=5.551115123e-23 pketa=-6.938893904e-30 dwg=0.0 dwb=0.0 pclm=6.151398981e-01 lpclm=-7.210786349e-8 pdiblc1=-2.150883798e-01 lpdiblc1=1.095415826e-07 wpdiblc1=1.110223025e-22 ppdiblc1=-8.326672685e-29 pdiblc2=-6.356604809e-03 lpdiblc2=2.826853610e-09 wpdiblc2=3.686287386e-24 ppdiblc2=-1.382357770e-30 pdiblcb=-8.794872769e-02 lpdiblcb=-2.938743745e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406427e+08 lpscbe1=1.198662602e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637210e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-8.497299977e-01 lkt1=8.486262334e-8 kt2=-4.272334130e-02 lkt2=2.651009219e-9 at=-3.181692162e+03 lat=6.108820679e-03 pat=7.275957614e-24 ute=-1.303565937e+00 lute=-2.963679149e-9 ua1=1.486947612e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 uc1=-1.025991505e-10 luc1=4.783040721e-17 wuc1=7.754818243e-32 puc1=3.877409121e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.106 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493649897e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810552122e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.754998478e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940225758e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372697511e-16 ags=1.250000000e+00 lags=2.938982391e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-08 pketa=-5.551115123e-29 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350075690e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301001387e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865618771e-18 drout=5.033266590e-01 ldrout=1.244684356e-16 pscbe1=7.914198799e+08 lpscbe1=1.229667664e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458478279e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407276948e-25 ub1=7.077531684e-19 lub1=1.999107579e-34 uc1=1.471862500e-10 luc1=-2.894304963e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.107 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-4.102081512e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.432828941e-07 wvth0=3.040372935e-06 pvth0=-3.693627463e-13 k1=0.90707349 k2=-1.995423928e+00 lk2=2.276604350e-07 wk2=1.141251635e-06 pk2=-1.386460961e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585356285e-01 ldsub=1.146481210e-11 wdsub=6.234481134e-11 pdsub=-7.574021750e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-7.534944890e-20 cit=0.0 voff='7.108895776e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.888433018e-07 wvoff=-4.613972220e-06 pvoff=5.605330291e-13 nfactor=2.603656528e+01 lnfactor=-2.771767059e-06 wnfactor=-1.334487157e-05 pnfactor=1.621215067e-12 eta0=1.342129091e-02 leta0=-1.630498760e-09 weta0=-8.866532836e-09 peta0=1.077159608e-15 etab=-0.043998 u0=2.851052724e-01 lu0=-3.101184626e-08 wu0=-1.573582368e-07 pu0=1.911682276e-14 ua=-1.847313362e-09 lua=8.348186473e-17 wua=3.721492690e-16 pua=-4.521092610e-23 ub=1.245014239e-18 lub=1.315444194e-25 wub=7.873095331e-25 pub=-9.564708593e-32 uc=2.775970619e-10 luc=-2.436924873e-17 wuc=-1.325181958e-16 puc=1.609910553e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.749294482e+05 lvsat=-1.008675050e-01 wvsat=-5.051463529e-01 pvsat=6.136820983e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=9.005330229e-06 lb0=-1.089573278e-12 wb0=-5.851253655e-12 pb0=7.108454016e-19 b1=3.247533933e-07 lb1=-3.945934784e-14 wb1=-2.146824738e-13 pb1=2.608091501e-20 keta=-2.700000006e-02 lketa=5.196704178e-18 dwg=0.0 dwb=0.0 pclm=-2.102611518e-01 lpclm=4.734419906e-08 wpclm=2.503586939e-07 ppclm=-3.041507629e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.141482776e-24 alpha1=0.85 beta0=1.390318599e+01 lbeta0=-4.865773908e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-1.201227025e+01 lkt1=1.408181014e-06 wkt1=7.274794410e-06 pkt1=-8.837856737e-13 kt2=-0.028878939 at=5.372048694e+04 lat=5.720299669e-12 ute=-8.308426021e-02 lute=-1.497528129e-07 wute=-8.077299354e-07 pute=9.812787893e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-4.801442190e-02 ltvoff=5.833080059e-09 wtvoff=3.027943091e-08 ptvoff=-3.678526944e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.108 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.109 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-7 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-8 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 uc=6.324132312e-11 luc=-2.932260536e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 b1=2.824547271e-08 lb1=-5.375173124e-14 wb1=-2.117582368e-28 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-7 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-7 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.110 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-7 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 uc=9.745036741e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-8 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=8.881784197e-22 ppclm=-1.421085472e-26 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116796e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 wuc1=2.067951531e-31 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.111 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 ub=1.752388505e-18 lub=-1.139532890e-24 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929613e-08 lb1=-3.422509015e-14 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-06 wpclm=7.105427358e-21 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-8 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-1 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 ub1=-1.471838908e-18 lub1=3.150583117e-24 wub1=6.162975822e-39 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-09 wtvoff=2.775557562e-23 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.112 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-8 k2=-7.388526331e-02 lk2=3.200507309e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-7 eta0=-1.412393437e-03 leta0=3.712885085e-09 peta0=6.938893904e-30 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=4.857225733e-23 petab=-3.122502257e-28 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-6 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=-1.110223025e-22 pketa=-2.775557562e-28 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-9 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=6.352747104e-27 palpha0=-7.199780052e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-08 wkt2=-4.440892099e-22 at=1.533204212e+05 lat=-8.532912747e-2 ute=-2.347817386e+00 lute=1.198707212e-6 ua1=-1.510649725e-09 lua1=2.628829754e-15 pua1=-6.617444900e-36 ub1=9.241642797e-19 lub1=-1.501223529e-24 wub1=-1.540743956e-39 pub1=-1.540743956e-45 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.113 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.724451032e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.919953230e-8 k1=6.241244142e-01 lk1=-6.584338284e-8 k2=-6.317640297e-02 lk2=2.192283100e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.340281270e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.282038687e-7 nfactor=-1.233075445e-02 lnfactor=2.173696432e-6 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=-9.159339953e-22 peta0=5.134781489e-28 etab=-1.583239050e-01 letab=6.962185878e-8 u0=2.995469753e-02 lu0=-2.435942066e-9 ua=-8.565838072e-10 lua=-2.614755107e-16 ub=1.909117804e-18 lub=1.054014256e-25 uc=2.808849156e-11 luc=1.079367420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.610106241e+04 lvsat=4.454635133e-2 a0=1.037003369e+00 la0=1.534590465e-7 ags=2.215750624e+00 lags=-9.092406921e-7 a1=0.0 a2=0.42385546 b0=4.720422506e-07 lb0=-2.084000450e-13 b1=2.945156506e-08 lb1=-1.300245365e-14 keta=-1.117400778e-01 lketa=4.619125186e-8 dwg=0.0 dwb=0.0 pclm=1.239890271e+00 lpclm=-3.479264068e-7 pdiblc1=6.380995512e-01 lpdiblc1=-2.671289443e-7 pdiblc2=8.798868558e-03 lpdiblc2=-3.864075705e-9 pdiblcb=8.317315893e-02 lpdiblcb=-7.848666098e-08 wpdiblcb=2.151057110e-22 ppdiblcb=1.283695372e-28 drout=8.488040648e-01 ldrout=6.675084449e-8 pscbe1=9.960958087e+08 lpscbe1=-2.468563664e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414640e-06 lalpha0=-1.346715357e-12 alpha1=0.85 beta0=1.697483351e+01 lbeta0=4.605433985e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=6.339107061e-02 lkt1=-3.182675446e-7 kt2=-1.865572788e-02 lkt2=-7.974505161e-9 at=1.086315090e+05 lat=-4.325514223e-2 ute=-8.665203951e-01 lute=-1.959131673e-7 ua1=1.678807431e-09 lua1=-3.739995058e-16 wua1=1.323488980e-29 ub1=-7.043401311e-19 lub1=3.199057494e-26 uc1=7.216247987e-11 luc1=-2.932440595e-17 kt1l=0.0 prt=0.0 tvoff=1.690720559e-03 ltvoff=-7.464294566e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.114 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.482941075e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.853720580e-8 k1=1.440277360e-01 lk1=1.461125792e-7 k2=7.969704024e-02 lk2=-4.115379395e-08 wk2=1.110223025e-22 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-1.169482067e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.178247696e-8 nfactor=5.439654304e+00 lnfactor=-2.332786435e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 petab=-6.938893904e-30 u0=2.047379937e-02 lu0=1.749741742e-9 ua=-1.652990168e-09 lua=9.012674784e-17 ub=2.069596195e-18 lub=3.455246251e-26 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.343617910e+05 lvsat=1.165615310e-3 a0=1.296210063e+00 la0=3.902291978e-8 ags=-6.815012482e-01 lags=3.698554480e-7 a1=0.0 a2=0.42385546 b0=1.286445378e-16 lb0=-2.463362796e-23 b1=-6.333203389e-18 lb1=1.212719784e-24 keta=5.112499917e-02 lketa=-2.571139952e-08 wketa=-1.665334537e-22 pketa=-6.938893904e-29 dwg=0.0 dwb=0.0 pclm=6.151398981e-01 lpclm=-7.210786349e-8 pdiblc1=-2.150883798e-01 lpdiblc1=1.095415826e-07 wpdiblc1=-4.440892099e-22 ppdiblc1=-3.330669074e-28 pdiblc2=-6.356604809e-03 lpdiblc2=2.826853610e-09 wpdiblc2=1.301042607e-23 ppdiblc2=1.951563910e-30 pdiblcb=-8.794872769e-02 lpdiblcb=-2.938743745e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406427e+08 lpscbe1=1.198662602e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637210e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-8.497299977e-01 lkt1=8.486262334e-08 wkt1=-7.105427358e-21 kt2=-4.272334130e-02 lkt2=2.651009219e-9 at=-3.181692162e+03 lat=6.108820679e-3 ute=-1.303565937e+00 lute=-2.963679149e-9 ua1=1.486947612e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 uc1=-1.025991505e-10 luc1=4.783040721e-17 wuc1=-3.618915180e-31 puc1=1.421716678e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.115 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493472261e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.812328479e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.755015826e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940225758e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372697511e-16 ags=1.250000000e+00 lags=2.939160026e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-8 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350031281e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301070776e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865618771e-18 drout=5.033266590e-01 ldrout=1.244675474e-16 pscbe1=7.914198799e+08 lpscbe1=1.229667664e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458478279e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407276172e-25 ub1=7.077531684e-19 lub1=1.999115282e-34 uc1=1.471862500e-10 luc1=-2.894718554e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.116 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.064529920e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.200487136e-08 wvth0=3.863364033e-07 pvth0=-4.693446430e-14 k1=0.90707349 k2=-1.526326585e-01 lk2=3.787094939e-09 wk2=-2.087150889e-08 pk2=2.535596129e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585349332e-01 ldsub=1.154929097e-11 wdsub=6.278333986e-11 pdsub=-7.627296826e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-7.534251001e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.871214957e-18 nfactor=4.840806852e-01 lnfactor=3.325020836e-07 wnfactor=2.769342895e-06 pnfactor=-3.364363909e-13 eta0=1.342125965e-02 leta0=-1.630495126e-09 weta0=-8.866513969e-09 peta0=1.077157316e-15 etab=-0.043998 u0=-1.155742062e-01 lu0=1.766510087e-08 wu0=9.532306408e-08 pu0=-1.158041776e-14 ua=9.033850581e-10 lua=-2.506894835e-16 wua=-1.362529177e-15 pua=1.655282196e-22 ub=-1.899937915e-18 lub=5.136120767e-25 wub=2.770616999e-24 pub=-3.365911768e-31 uc=2.790688779e-10 luc=-2.454805377e-17 wuc=-1.334463700e-16 puc=1.621186571e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.562698740e+05 lvsat=-1.356042801e-02 wvsat=-5.193662834e-02 pvsat=6.309573230e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=9.005212994e-06 lb0=-1.089559035e-12 wb0=-5.851179724e-12 pb0=7.108364199e-19 b1=3.247540737e-07 lb1=-3.945943049e-14 wb1=-2.146829028e-13 pb1=2.608096713e-20 keta=-2.700000006e-02 lketa=5.196731934e-18 dwg=0.0 dwb=0.0 pclm=-2.102611435e-01 lpclm=4.734419805e-08 wpclm=2.503586887e-07 ppclm=-3.041507566e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.141588655e-24 alpha1=0.85 beta0=1.390318599e+01 lbeta0=-4.865773908e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.177049964e+00 lkt1=2.133394424e-07 wkt1=1.072389772e-06 pkt1=-1.302803438e-13 kt2=-0.028878939 at=5.372048694e+04 lat=5.720416084e-12 ute=-7.411315990e-02 lute=-1.508426760e-07 wute=-8.133873983e-07 pute=9.881518147e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.117 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.118 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-7 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-8 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 uc=6.324132312e-11 luc=-2.932260536e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 b1=2.824547271e-08 lb1=-5.375173124e-14 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-7 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+03 ppscbe1=7.629394531e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-07 wkt2=-1.110223025e-22 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.119 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-07 pk2=-4.440892099e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-7 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 uc=9.745036742e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-8 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=-4.440892099e-22 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116797e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.120 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 ub=1.752388505e-18 lub=-1.139532890e-24 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929613e-08 lb1=-3.422509015e-14 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-6 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-08 wpdiblcb=1.110223025e-22 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-1 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 ub1=-1.471838908e-18 lub1=3.150583117e-24 pub1=6.162975822e-45 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.121 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-8 k2=-7.388526331e-02 lk2=3.200507309e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-7 eta0=-1.412393437e-03 leta0=3.712885085e-09 peta0=-6.938893904e-30 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=-2.775557562e-23 petab=-6.938893904e-30 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 pua=-1.654361225e-36 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-6 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=8.326672685e-23 pketa=2.220446049e-28 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-9 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=4.658681210e-27 palpha0=-3.388131789e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-8 at=1.533204212e+05 lat=-8.532912747e-2 ute=-2.347817386e+00 lute=1.198707212e-06 wute=7.105427358e-21 ua1=-1.510649725e-09 lua1=2.628829754e-15 pua1=-1.654361225e-36 ub1=9.241642797e-19 lub1=-1.501223529e-24 wub1=7.703719778e-40 pub1=3.081487911e-45 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.122 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.700669189e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.091406714e-06 wvth0=-7.002119710e-07 pvth0=6.592397678e-13 k1=6.241244150e-01 lk1=-6.584338359e-08 wk1=-4.894573635e-16 pk1=4.608171622e-22 k2=-6.551785979e-02 lk2=2.412727982e-08 wk2=1.453183031e-09 pk2=-1.368151479e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802130e-01 ldsub=4.182060754e-08 wdsub=-1.443645203e-16 pdsub=1.359161672e-22 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-5.046405876e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.470692946e-06 wvoff=2.862589227e-06 pvoff=-2.695087681e-12 nfactor=-7.114487967e+01 lnfactor=6.914399538e-05 wnfactor=4.414713610e-05 pnfactor=-4.156391058e-11 eta0=-4.278900077e-01 leta0=4.052355882e-07 weta0=3.302971369e-16 peta0=-3.109717345e-22 etab=-1.583239051e-01 letab=6.962185888e-08 wetab=6.636380334e-17 petab=-6.248068729e-23 u0=-1.511767842e-02 lu0=3.999906888e-08 wu0=2.797335883e-08 pu0=-2.633652571e-14 ua=-5.622285063e-10 lua=-5.386069054e-16 wua=-1.826863191e-16 pua=1.719966118e-22 ub=1.641290178e-18 lub=3.575573857e-25 wub=1.662223951e-25 pub=-1.564960578e-31 uc=2.808849168e-11 luc=1.079367408e-17 wuc=-7.439703788e-26 puc=7.004379311e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-7.346743722e+04 lvsat=1.477035598e-01 wvsat=6.800171706e-02 pvsat=-6.402266459e-8 a0=1.037003363e+00 la0=1.534590520e-07 wa0=3.598238152e-15 pa0=-3.387683023e-21 ags=2.215750599e+00 lags=-9.092406680e-07 wags=1.589961585e-14 pags=-1.496926672e-20 a1=0.0 a2=0.42385546 b0=4.720422487e-07 lb0=-2.084000432e-13 wb0=1.198875187e-21 pb0=-1.128723918e-27 b1=2.945156515e-08 lb1=-1.300245374e-14 wb1=-5.902093813e-23 pb1=5.556737304e-29 keta=-1.117400787e-01 lketa=4.619125269e-08 wketa=5.486051613e-16 pketa=-5.165042838e-22 dwg=0.0 dwb=0.0 pclm=1.239890278e+00 lpclm=-3.479264132e-07 wpclm=-4.203020154e-15 ppclm=3.957087102e-21 pdiblc1=6.380995499e-01 lpdiblc1=-2.671289431e-07 wpdiblc1=7.878195873e-16 ppdiblc1=-7.417204628e-22 pdiblc2=8.798868589e-03 lpdiblc2=-3.864075734e-09 wpdiblc2=-1.898578517e-17 ppdiblc2=1.787485437e-23 pdiblcb=8.317315868e-02 lpdiblcb=-7.848666075e-08 wpdiblcb=1.525364756e-16 ppdiblcb=-1.436108199e-22 drout=8.488040656e-01 ldrout=6.675084369e-08 wdrout=-5.294680250e-16 pdrout=4.984848090e-22 pscbe1=9.960957989e+08 lpscbe1=-2.468563571e+02 wpscbe1=6.096603394e-06 ppscbe1=-5.739866257e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414628e-06 lalpha0=-1.346715347e-12 walpha0=7.156140914e-21 palpha0=-6.737422035e-27 alpha1=0.85 beta0=1.697483357e+01 lbeta0=4.605433502e-07 wbeta0=-3.186312370e-14 pbeta0=2.999860271e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=1.010169003e+01 lkt1=-9.769185478e-06 wkt1=-6.230089559e-06 pkt1=5.865542099e-12 kt2=-1.865572789e-02 lkt2=-7.974505148e-09 wkt2=8.334000157e-18 pkt2=-7.846279182e-24 at=1.086315079e+05 lat=-4.325514127e-02 wat=6.332173944e-10 pat=-5.961654242e-16 ute=-8.665203930e-01 lute=-1.959131693e-07 wute=-1.308855246e-15 pute=1.232269398e-21 ua1=1.678807427e-09 lua1=-3.739995017e-16 wua1=2.711511283e-24 pua1=-2.552851424e-30 ub1=-7.043401320e-19 lub1=3.199057584e-26 wub1=5.949028116e-34 pub1=-5.600912427e-40 uc1=7.216247998e-11 luc1=-2.932440605e-17 wuc1=-6.588824451e-26 puc1=6.203285907e-32 kt1l=0.0 prt=0.0 tvoff=3.561664957e-02 ltvoff=-3.268721666e-08 wtvoff=-2.105551718e-08 ptvoff=1.982347464e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.123 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-1.708154065e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.135410289e-07 wvth0=1.400423942e-06 pvth0=-2.681615790e-13 k1=1.440277344e-01 lk1=1.461125795e-07 wk1=9.789147271e-16 pk1=-1.874487232e-22 k2=8.437995389e-02 lk2=-4.205050635e-08 wk2=-2.906366061e-09 pk2=5.565284116e-16 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001172e-01 ldsub=5.015590555e-08 wdsub=2.887272643e-16 pdsub=-5.528710822e-23 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='9.107807290e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.778194008e-06 wvoff=-5.725178454e-06 pvoff=1.096291521e-12 nfactor=1.477047521e+02 lnfactor=-2.747505317e-05 wnfactor=-8.829427220e-05 pnfactor=1.690711701e-11 eta0=8.647808887e-01 leta0=-1.654605151e-07 weta0=-6.605986869e-16 peta0=1.264952587e-22 etab=3.259628934e-02 letab=-1.466673409e-08 wetab=-1.327278842e-16 petab=2.541552819e-23 u0=1.106185513e-01 lu0=-1.551171622e-08 wu0=-5.594671766e-08 pu0=1.071301318e-14 ua=-2.241700769e-09 lua=2.028565861e-16 wua=3.653726382e-16 pua=-6.996374499e-23 ub=2.605251447e-18 lub=-6.801801901e-26 wub=-3.324447901e-25 pub=6.365852308e-32 uc=2.188162303e-11 luc=1.353391970e-17 wuc=1.487942826e-25 puc=-2.849197771e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.534987903e+05 lvsat=-4.079605213e-02 wvsat=-1.360034341e-01 pvsat=2.604275359e-8 a0=1.296210075e+00 la0=3.902291756e-08 wa0=-7.196469198e-15 pa0=1.378023029e-21 ags=-6.815011970e-01 lags=3.698554382e-07 wags=-3.179922814e-14 pags=6.089106663e-21 a1=0.0 a2=0.42385546 b0=3.992045838e-15 lb0=-7.644208893e-22 wb0=-2.397750476e-21 pb0=4.591356476e-28 b1=-1.965294343e-16 lb1=3.763263525e-23 wb1=1.180418672e-22 pb1=-2.260336498e-29 keta=5.112500094e-02 lketa=-2.571139986e-08 wketa=-1.097210628e-15 pketa=2.101004787e-22 dwg=0.0 dwb=0.0 pclm=6.151398845e-01 lpclm=-7.210786090e-08 wpclm=8.406045637e-15 ppclm=-1.609639977e-21 pdiblc1=-2.150883772e-01 lpdiblc1=1.095415821e-07 wpdiblc1=-1.575638287e-15 ppdiblc1=3.017127936e-22 pdiblc2=-6.356604870e-03 lpdiblc2=2.826853621e-09 wpdiblc2=3.797156166e-17 ppdiblc2=-7.271020429e-24 pdiblcb=-8.794872720e-02 lpdiblcb=-2.938743839e-09 wpdiblcb=-3.050728559e-16 ppdiblcb=5.841716000e-23 drout=1.380423787e+00 ldrout=-1.679518205e-07 wdrout=1.058936050e-15 pdrout=-2.027702450e-22 pscbe1=1.654406624e+08 lpscbe1=1.198662565e+02 wpscbe1=-1.219320869e-05 ppscbe1=2.334828854e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637233e-06 lalpha0=-1.311494744e-12 walpha0=-1.431230893e-20 palpha0=2.740605594e-27 alpha1=0.85 beta0=2.085046081e+01 lbeta0=-1.250491818e-06 wbeta0=6.372613370e-14 pbeta0=-1.220266199e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.092632791e+01 lkt1=3.929250052e-06 wkt1=1.246017912e-05 pkt1=-2.385949859e-12 kt2=-4.272334128e-02 lkt2=2.651009214e-09 wkt2=-1.666800031e-17 pkt2=3.191696907e-24 at=-3.181690121e+03 lat=6.108820288e-03 wat=-1.266434905e-09 pat=2.425045532e-16 ute=-1.303565941e+00 lute=-2.963678342e-09 wute=2.617710493e-15 pute=-5.012541493e-22 ua1=1.486947620e-09 lua1=-2.892960831e-16 wua1=-5.423022566e-24 pua1=1.038432615e-30 ub1=-1.657962220e-18 lub1=4.530013771e-25 wub1=-1.189796379e-33 pub1=2.278313494e-40 uc1=-1.025991507e-10 luc1=4.783040725e-17 wuc1=1.317766441e-25 puc1=-2.523332553e-32 kt1l=0.0 prt=0.0 tvoff=-6.785185803e-02 ltvoff=1.299268089e-08 wtvoff=4.211103435e-08 ptvoff=-8.063673524e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.124 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493472261e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810552122e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.754981131e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940225758e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372715275e-16 ags=1.250000000e+00 lags=2.938982391e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-8 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350031281e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.300931998e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865618771e-18 drout=5.033266590e-01 ldrout=1.244684356e-16 pscbe1=7.914198799e+08 lpscbe1=1.229572296e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458478279e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407276689e-25 ub1=7.077531684e-19 lub1=1.999099875e-34 uc1=1.471862500e-10 luc1=-2.894511758e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.125 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-7.950669847e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.459637032e-08 wvth0=5.017489380e-07 pvth0=-6.095547148e-14 k1=0.90707349 k2=-4.050020702e-01 lk2=3.444644529e-08 wk2=1.357570239e-07 pk2=-1.649257780e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585343557e-01 ldsub=1.161944248e-11 wdsub=6.314172084e-11 pdsub=-7.670835098e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-7.534944890e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.870770867e-18 nfactor=1.742783651e+01 lnfactor=-1.725927036e-06 wnfactor=-7.746494169e-06 pnfactor=9.410905906e-13 eta0=1.342126029e-02 leta0=-1.630495203e-09 weta0=-8.866514362e-09 peta0=1.077157364e-15 etab=-0.043998 u0=1.262843539e-01 lu0=-1.171732816e-08 wu0=-5.478209779e-08 pu0=6.655257932e-15 ua=9.033804188e-10 lua=-2.506889199e-16 wua=-1.362526298e-15 pua=1.655278698e-22 ub=-1.899821614e-18 lub=5.135979478e-25 wub=2.770544819e-24 pub=-3.365824079e-31 uc=2.802962414e-10 luc=-2.469716124e-17 wuc=-1.342081111e-16 puc=1.630440658e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.138312164e+05 lvsat=-2.055332526e-02 wvsat=-8.766103941e-02 pvsat=1.064958903e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=9.005291601e-06 lb0=-1.089568585e-12 wb0=-5.851228510e-12 pb0=7.108423467e-19 b1=3.247514418e-07 lb1=-3.945911075e-14 wb1=-2.146812694e-13 pb1=2.608076869e-20 keta=-2.700000006e-02 lketa=5.196676423e-18 dwg=0.0 dwb=0.0 pclm=-2.102611471e-01 lpclm=4.734419849e-08 wpclm=2.503586909e-07 ppclm=-3.041507593e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.141482776e-24 alpha1=0.85 beta0=1.390318599e+01 lbeta0=-4.865773908e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=3.106190437e+00 lkt1=-4.285003010e-07 wkt1=-2.206558285e-06 pkt1=2.680659398e-13 kt2=-0.028878939 at=5.372048694e+04 lat=5.720299669e-12 ute=-6.663208752e-02 lute=-1.517515215e-07 wute=-8.180303912e-07 pute=9.937924011e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.126 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.127 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-7 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-08 wu0=-5.551115123e-23 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 uc=6.324132312e-11 luc=-2.932260536e-16 wuc=1.033975766e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 b1=2.824547271e-08 lb1=-5.375173124e-14 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-7 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+03 ppscbe1=3.814697266e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-7 at=1.981626675e+05 lat=-4.618980097e-01 wat=4.656612873e-16 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 wuc1=1.033975766e-31 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.128 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-07 pk2=-2.220446049e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-07 wvoff=8.881784197e-22 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 uc=9.745036741e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-8 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=2.220446049e-22 ppclm=4.440892099e-27 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-08 ppdiblc2=2.775557562e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116796e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 wua1=-3.308722450e-30 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 wuc1=5.169878828e-32 puc1=2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.129 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-06 wdsub=1.776356839e-21 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 ub=1.752388505e-18 lub=-1.139532890e-24 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929614e-08 lb1=-3.422509015e-14 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-6 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-8 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-1 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 ub1=-1.471838908e-18 lub1=3.150583117e-24 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-09 wtvoff=-6.938893904e-24 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.130 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-8 k2=-7.388526331e-02 lk2=3.200507309e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-07 wnfactor=7.105427358e-21 eta0=-1.412393438e-03 leta0=3.712885085e-09 weta0=-1.734723476e-24 peta0=-3.469446952e-30 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=3.642919300e-23 petab=1.075528555e-28 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-6 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=1.387778781e-23 pketa=9.714451465e-29 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-9 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=-1.058791184e-27 palpha0=3.176373552e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-8 at=1.533204212e+05 lat=-8.532912747e-2 ute=-2.347817386e+00 lute=1.198707212e-6 ua1=-1.510649725e-09 lua1=2.628829754e-15 wua1=-1.654361225e-30 pua1=2.067951531e-36 ub1=9.241642797e-19 lub1=-1.501223529e-24 wub1=-3.851859889e-40 pub1=7.703719778e-46 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.131 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.348772052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.170117734e-9 k1=6.241244142e-01 lk1=-6.584338282e-8 k2=-6.309843653e-02 lk2=2.184942669e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.804439774e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.639345798e-8 nfactor=2.356259295e+00 lnfactor=-5.629793918e-8 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=-4.093947403e-22 peta0=-2.983724379e-28 etab=-1.583239050e-01 letab=6.962185877e-8 u0=3.145552919e-02 lu0=-3.848954058e-9 ua=-8.663853263e-10 lua=-2.522475177e-16 ub=1.918035997e-18 lub=9.700507105e-26 uc=2.808849155e-11 luc=1.079367420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.974950271e+04 lvsat=4.111139587e-2 a0=1.037003369e+00 la0=1.534590463e-7 ags=2.215750625e+00 lags=-9.092406929e-7 a1=0.0 a2=0.42385546 b0=4.720422507e-07 lb0=-2.084000451e-13 b1=2.945156505e-08 lb1=-1.300245365e-14 keta=-1.117400778e-01 lketa=4.619125183e-8 dwg=0.0 dwb=0.0 pclm=1.239890271e+00 lpclm=-3.479264066e-7 pdiblc1=6.380995512e-01 lpdiblc1=-2.671289443e-7 pdiblc2=8.798868557e-03 lpdiblc2=-3.864075704e-9 pdiblcb=8.317315894e-02 lpdiblcb=-7.848666099e-08 wpdiblcb=-3.816391647e-23 ppdiblcb=-4.813857646e-29 drout=8.488040648e-01 ldrout=6.675084452e-8 pscbe1=9.960958090e+08 lpscbe1=-2.468563667e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414640e-06 lalpha0=-1.346715358e-12 walpha0=-1.355252716e-26 alpha1=0.85 beta0=1.697483351e+01 lbeta0=4.605434001e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.708668097e-01 lkt1=-3.568429924e-9 kt2=-1.865572788e-02 lkt2=-7.974505161e-9 at=1.086315090e+05 lat=-4.325514226e-2 ute=-8.665203951e-01 lute=-1.959131673e-7 ua1=1.678807431e-09 lua1=-3.739995059e-16 ub1=-7.043401311e-19 lub1=3.199057490e-26 uc1=7.216247987e-11 luc1=-2.932440595e-17 kt1l=0.0 prt=0.0 tvoff=5.610461820e-04 ltvoff=3.171431537e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.132 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.234299035e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.292465884e-8 k1=1.440277361e-01 lk1=1.461125792e-7 k2=7.954110737e-02 lk2=-4.112393499e-08 pk2=2.081668171e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-4.241165060e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.703595200e-8 nfactor=7.024742053e-01 lnfactor=6.738250248e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 wetab=-6.938893904e-24 petab=8.673617380e-30 u0=1.747213606e-02 lu0=2.324518243e-9 ua=-1.633387130e-09 lua=8.637304047e-17 ub=2.051759808e-18 lub=3.796788098e-26 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.270649104e+05 lvsat=2.562865788e-3 a0=1.296210063e+00 la0=3.902291985e-8 ags=-6.815012499e-01 lags=3.698554483e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.112499912e-02 lketa=-2.571139951e-08 wketa=5.551115123e-23 pketa=2.081668171e-29 dwg=0.0 dwb=0.0 pclm=6.151398985e-01 lpclm=-7.210786358e-8 pdiblc1=-2.150883799e-01 lpdiblc1=1.095415826e-07 wpdiblc1=-1.110223025e-22 ppdiblc1=8.326672685e-29 pdiblc2=-6.356604807e-03 lpdiblc2=2.826853609e-09 wpdiblc2=-2.927345866e-24 ppdiblc2=-4.878909776e-31 pdiblcb=-8.794872771e-02 lpdiblcb=-2.938743742e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406421e+08 lpscbe1=1.198662603e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637209e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-1.812142371e-01 lkt1=-4.314878560e-8 kt2=-4.272334130e-02 lkt2=2.651009219e-9 at=-3.181692230e+03 lat=6.108820692e-3 ute=-1.303565937e+00 lute=-2.963679176e-9 ua1=1.486947611e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 wub1=-1.540743956e-39 pub1=3.851859889e-46 uc1=-1.025991505e-10 luc1=4.783040720e-17 wuc1=3.877409121e-32 puc1=1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=2.259348754e-03 ltvoff=-4.326336554e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.133 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493649897e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810108033e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.754998478e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940281269e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372715275e-16 ags=1.250000000e+00 lags=2.938982391e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-8 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350031281e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301001387e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865729793e-18 drout=5.033266590e-01 ldrout=1.244684356e-16 pscbe1=7.914198799e+08 lpscbe1=1.229667664e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458478279e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407276948e-25 ub1=7.077531684e-19 lub1=1.999099875e-34 uc1=1.471862500e-10 luc1=-2.894511758e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.134 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='2.546308249e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.644033844e-07 wvth0=-1.075399546e-06 pvth0=1.306459892e-13 k1=0.90707349 k2=1.170170090e+00 lk2=-1.569149197e-07 wk2=-8.103417809e-07 pk2=9.844518159e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585332767e-01 ldsub=1.175052483e-11 wdsub=6.378979761e-11 pdsub=-7.749567353e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-7.534771418e-20 cit=0.0 voff='-5.826104817e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.825781802e-07 wvoff=3.374695829e-06 pvoff=-4.099782975e-13 nfactor=-5.107157664e+01 lnfactor=6.595792669e-06 wnfactor=3.339644535e-05 pnfactor=-4.057200559e-12 eta0=1.342123430e-02 leta0=-1.630492045e-09 weta0=-8.866498752e-09 peta0=1.077155467e-15 etab=-0.043998 u0=-3.304309512e-01 lu0=4.376718740e-08 wu0=2.195357294e-07 pu0=-2.667051762e-14 ua=4.454467095e-09 lua=-6.820962359e-16 wua=-3.495422590e-15 pua=4.246449088e-22 ub=-6.836087032e-18 lub=1.113285088e-24 wub=5.735423790e-24 pub=-6.967736945e-31 uc=2.825842743e-10 luc=-2.497512520e-17 wuc=-1.355823768e-16 puc=1.647136063e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.760033047e+05 lvsat=7.540051138e-02 wvsat=3.867388487e-01 pvsat=-4.698335577e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=9.005334457e-06 lb0=-1.089573791e-12 wb0=-5.851254250e-12 pb0=7.108454738e-19 b1=3.247549466e-07 lb1=-3.945953653e-14 wb1=-2.146833744e-13 pb1=2.608102443e-20 keta=-2.700000006e-02 lketa=5.196704178e-18 dwg=0.0 dwb=0.0 pclm=-2.102611534e-01 lpclm=4.734419925e-08 wpclm=2.503586947e-07 ppclm=-3.041507638e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.141482776e-24 alpha1=0.85 beta0=1.390318599e+01 lbeta0=-4.865773908e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=7.085908648e+00 lkt1=-9.119803476e-07 wkt1=-4.596904393e-06 pkt1=5.584595271e-13 kt2=-0.028878939 at=5.372048694e+04 lat=5.720299669e-12 ute=-5.268595525e-02 lute=-1.534457813e-07 wute=-8.264068846e-07 pute=1.003968668e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=2.492665059e-02 ltvoff=-3.028239073e-09 wtvoff=-1.497174400e-08 ptvoff=1.818857291e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.135 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.136 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-7 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-8 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 uc=6.324132312e-11 luc=-2.932260536e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 b1=2.824547271e-08 lb1=-5.375173124e-14 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-07 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+03 ppscbe1=-1.525878906e-17 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-7 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 wuc1=2.067951531e-31 puc1=-1.654361225e-36 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.137 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-7 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 wub=1.232595164e-38 uc=9.745036741e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-8 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=-4.440892099e-22 ppclm=-7.105427358e-27 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116797e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.138 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 ub=1.752388505e-18 lub=-1.139532890e-24 wub=1.232595164e-38 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929613e-08 lb1=-3.422509015e-14 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-6 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-8 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-1 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 ub1=-1.471838908e-18 lub1=3.150583117e-24 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.139 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-8 k2=-7.388526331e-02 lk2=3.200507309e-08 wk2=-4.440892099e-22 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-7 eta0=-1.412393438e-03 leta0=3.712885085e-09 peta0=-3.469446952e-30 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=1.318389842e-22 petab=-1.075528555e-28 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-06 pags=-3.552713679e-27 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=5.551115123e-23 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-9 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=-8.470329473e-28 palpha0=-9.740878893e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-8 at=1.533204212e+05 lat=-8.532912747e-02 wat=9.313225746e-16 ute=-2.347817386e+00 lute=1.198707212e-6 ua1=-1.510649725e-09 lua1=2.628829754e-15 wua1=3.308722450e-30 pua1=6.617444900e-36 ub1=9.241642797e-19 lub1=-1.501223529e-24 wub1=-1.540743956e-39 pub1=-1.540743956e-45 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.140 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.348772052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.170117734e-9 k1=6.241244142e-01 lk1=-6.584338282e-8 k2=-6.309843653e-02 lk2=2.184942669e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.804439774e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.639345798e-8 nfactor=2.356259295e+00 lnfactor=-5.629793918e-8 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=3.330669074e-22 peta0=3.053113318e-28 etab=-1.583239050e-01 letab=6.962185877e-8 u0=3.145552919e-02 lu0=-3.848954058e-9 ua=-8.663853263e-10 lua=-2.522475177e-16 ub=1.918035997e-18 lub=9.700507105e-26 uc=2.808849155e-11 luc=1.079367420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.974950271e+04 lvsat=4.111139587e-2 a0=1.037003369e+00 la0=1.534590463e-7 ags=2.215750625e+00 lags=-9.092406929e-7 a1=0.0 a2=0.42385546 b0=4.720422507e-07 lb0=-2.084000451e-13 b1=2.945156505e-08 lb1=-1.300245365e-14 keta=-1.117400778e-01 lketa=4.619125183e-8 dwg=0.0 dwb=0.0 pclm=1.239890271e+00 lpclm=-3.479264066e-7 pdiblc1=6.380995512e-01 lpdiblc1=-2.671289443e-7 pdiblc2=8.798868557e-03 lpdiblc2=-3.864075704e-9 pdiblcb=8.317315894e-02 lpdiblcb=-7.848666099e-08 wpdiblcb=1.283695372e-22 ppdiblcb=-1.708702624e-28 drout=8.488040648e-01 ldrout=6.675084452e-8 pscbe1=9.960958090e+08 lpscbe1=-2.468563667e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414640e-06 lalpha0=-1.346715358e-12 alpha1=0.85 beta0=1.697483351e+01 lbeta0=4.605434001e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.708668097e-01 lkt1=-3.568429924e-9 kt2=-1.865572788e-02 lkt2=-7.974505161e-9 at=1.086315090e+05 lat=-4.325514226e-2 ute=-8.665203951e-01 lute=-1.959131673e-7 ua1=1.678807431e-09 lua1=-3.739995059e-16 ub1=-7.043401311e-19 lub1=3.199057490e-26 uc1=7.216247987e-11 luc1=-2.932440595e-17 kt1l=0.0 prt=0.0 tvoff=5.610461820e-04 ltvoff=3.171431537e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.141 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.234299035e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.292465884e-8 k1=1.440277361e-01 lk1=1.461125792e-7 k2=7.954110737e-02 lk2=-4.112393499e-08 wk2=1.110223025e-22 pk2=-5.551115123e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-09 pcdscd=6.938893904e-30 cit=0.0 voff='-4.241165060e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.703595200e-8 nfactor=7.024742053e-01 lnfactor=6.738250248e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 wetab=2.081668171e-23 petab=1.994931997e-29 u0=1.747213606e-02 lu0=2.324518243e-9 ua=-1.633387130e-09 lua=8.637304047e-17 ub=2.051759808e-18 lub=3.796788098e-26 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.270649104e+05 lvsat=2.562865788e-3 a0=1.296210063e+00 la0=3.902291985e-8 ags=-6.815012499e-01 lags=3.698554483e-07 wags=-1.776356839e-21 pags=-4.440892099e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.112499912e-02 lketa=-2.571139951e-08 wketa=5.551115123e-23 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=6.151398985e-01 lpclm=-7.210786358e-08 wpclm=-3.552713679e-21 pdiblc1=-2.150883799e-01 lpdiblc1=1.095415826e-07 wpdiblc1=4.440892099e-22 ppdiblc1=1.665334537e-28 pdiblc2=-6.356604807e-03 lpdiblc2=2.826853609e-09 wpdiblc2=4.770489559e-24 ppdiblc2=-5.746271514e-30 pdiblcb=-8.794872771e-02 lpdiblcb=-2.938743742e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406421e+08 lpscbe1=1.198662603e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637209e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-1.812142371e-01 lkt1=-4.314878560e-8 kt2=-4.272334130e-02 lkt2=2.651009219e-9 at=-3.181692230e+03 lat=6.108820692e-3 ute=-1.303565937e+00 lute=-2.963679176e-9 ua1=1.486947611e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 pub1=7.703719778e-46 uc1=-1.025991505e-10 luc1=4.783040720e-17 wuc1=-1.550963649e-31 puc1=-3.877409121e-38 kt1l=0.0 prt=0.0 tvoff=2.259348754e-03 ltvoff=-4.326336554e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.142 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493472261e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810552122e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.754946437e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940225758e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372697511e-16 ags=1.250000000e+00 lags=2.939160026e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-8 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350031281e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.300793221e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865618771e-18 drout=5.033266590e-01 ldrout=1.244693237e-16 pscbe1=7.914198799e+08 lpscbe1=1.229476929e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.458478279e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407277206e-25 ub1=7.077531684e-19 lub1=1.999099875e-34 uc1=1.471862500e-10 luc1=-2.895132144e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.143 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-6.958188337e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.902598879e-07 wvth0=4.348170351e-06 pvth0=-5.282418232e-13 k1=0.90707349 k2=-4.256628991e+00 lk2=5.023651935e-07 wk2=2.286363432e-06 pk2=-2.777611479e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.104959957e+00 ldsub=-2.000060412e-07 wdsub=-9.394399597e-07 pdsub=1.141288029e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-7.535638780e-20 cit=0.0 voff='1.664819445e+01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.047734540e-06 wvoff=-9.449858509e-06 pvoff=1.148025511e-12 nfactor=1.762249807e+02 lnfactor=-2.101755690e-05 wnfactor=-9.630624376e-05 pnfactor=1.169986033e-11 eta0=-9.291588981e-03 leta0=1.128798003e-09 weta0=4.094165021e-09 peta0=-4.973837317e-16 etab=-0.043998 u0=1.129870254e+00 lu0=-1.336389649e-07 wu0=-6.137588681e-07 pu0=7.456310986e-14 ua=-1.337283455e-08 lua=1.483671332e-15 wua=6.677406203e-15 pua=-8.112113700e-22 ub=2.624088074e-17 lub=-2.905103418e-24 wub=-1.313935248e-23 pub=1.596247376e-30 uc=-1.469740513e-10 luc=2.721019754e-17 wuc=1.095373496e-16 puc=-1.330725445e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.569057000e+06 lvsat=-2.945316849e-01 wvsat=-1.350870003e+00 pvsat=1.641117932e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-8.567905533e-06 lb0=1.045328842e-12 wb0=4.176598832e-12 pb0=-5.073982857e-19 b1=1.086901143e-08 lb1=-1.326789817e-15 wb1=-3.557001551e-14 pb1=4.321258904e-21 keta=-7.029949672e-01 lketa=8.212392458e-08 wketa=3.857443601e-07 pketa=-4.686253933e-14 dwg=0.0 dwb=0.0 pclm=2.588624598e-02 lpclm=1.865559629e-08 wpclm=1.156054319e-07 ppclm=-1.404444150e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.999998012e-08 lalpha0=2.415482691e-21 walpha0=1.135112749e-20 palpha0=-1.379003043e-27 alpha1=0.85 beta0=1.390318580e+01 lbeta0=-4.865750820e-09 wbeta0=1.084465566e-13 pbeta0=-1.317474130e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.267582301e+01 lkt1=2.703653385e-06 wkt1=1.238609207e-05 pkt1=-1.504736781e-12 kt2=-0.028878939 at=5.372048908e+04 lat=-2.546512987e-10 wat=-1.222989522e-09 pat=1.485762186e-16 ute=-1.141949138e+00 lute=-2.111555432e-08 wute=-2.048384560e-07 pute=2.488500467e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-7.477995176e-02 ltvoff=9.084717220e-09 wtvoff=4.192403392e-08 ptvoff=-5.093183184e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.144 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.145 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.941722858e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.600512189e-7 k1=6.121394710e-01 lk1=-8.800526942e-7 k2=-6.142183918e-02 lk2=3.446086836e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.219088418e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.236172364e-7 nfactor=2.751881615e+00 lnfactor=-1.489951008e-7 eta0=0.08 etab=-0.07 u0=2.447623674e-02 lu0=3.311808729e-8 ua=-1.241716814e-09 lua=3.742273392e-15 ub=1.952403039e-18 lub=-2.382469934e-24 wub=6.162975822e-39 uc=6.324132312e-11 luc=-2.932260536e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390792275e+00 la0=-5.621958632e-7 ags=3.209695092e-01 lags=4.768107168e-7 a1=0.0 a2=0.42385546 b0=7.046139034e-08 lb0=3.353379550e-14 b1=2.824547271e-08 lb1=-5.375173124e-14 keta=-2.668570919e-03 lketa=-3.745069062e-8 dwg=0.0 dwb=0.0 pclm=-9.596620000e-03 lpclm=5.278834396e-07 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=5.534321625e-04 lpdiblc2=8.114096878e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.280520219e+07 lpscbe1=5.938678270e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832298772e-01 lkt1=-6.281812932e-8 kt2=-3.543871383e-02 lkt2=1.180692079e-7 at=1.981626675e+05 lat=-4.618980097e-1 ute=-1.016329962e+00 lute=-1.975603773e-6 ua1=1.030268522e-09 lua1=1.809320489e-15 wua1=3.308722450e-30 ub1=-3.834803979e-19 lub1=-3.708909047e-24 uc1=6.915598073e-11 luc1=-7.046846291e-16 kt1l=0.0 prt=0.0 tvoff=1.685329285e-03 ltvoff=1.812223848e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.146 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.204864831e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.107738936e-8 k1=4.375091496e-01 lk1=5.067715585e-7 k2=9.832922552e-03 lk2=-2.212600092e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.561695447e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.484636565e-7 nfactor=2.921710646e+00 lnfactor=-1.497689971e-6 eta0=0.08 etab=-0.07 u0=2.728047949e-02 lu0=1.084823276e-8 ua=-9.755391182e-10 lua=1.628426944e-15 ub=1.838757400e-18 lub=-1.479954680e-24 uc=9.745036741e-12 luc=1.316139557e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408683435e+00 la0=-7.042782575e-7 ags=3.611449106e-01 lags=1.577583297e-7 a1=0.0 a2=0.42385546 b0=3.887954118e-08 lb0=2.843406085e-13 b1=1.348386815e-10 lb1=1.694884753e-13 keta=-1.737606701e-02 lketa=7.934868368e-8 dwg=0.0 dwb=0.0 pclm=-6.880116586e-01 lpclm=5.915506971e-06 wpclm=2.220446049e-22 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.615309433e-03 lpdiblc2=2.533712789e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.393250764e+08 lpscbe1=2.833056325e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.863116796e-01 lkt1=-3.834403846e-8 kt2=-9.889062257e-03 lkt2=-8.483299237e-8 at=140000.0 ute=-1.231301758e+00 lute=-2.684082692e-7 ua1=1.513656099e-09 lua1=-2.029495179e-15 ub1=-1.025915981e-18 lub1=1.392984140e-24 uc1=-7.075299815e-11 luc1=4.064005679e-16 kt1l=0.0 prt=0.0 tvoff=5.800682213e-03 ltvoff=-1.455977918e-08 wtvoff=-1.387778781e-23 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.147 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.295229188e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.546040489e-8 k1=5.592721859e-01 lk1=2.684425528e-8 k2=-3.553077567e-02 lk2=-4.245962771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.512229000e-01 ldsub=-1.147850983e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.486482770e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.188186849e-7 nfactor=2.345173169e+00 lnfactor=7.747244207e-7 eta0=1.571740685e-01 leta0=-3.041805106e-7 etab=-1.374666385e-01 letab=2.659188111e-7 u0=2.976419541e-02 lu0=1.058701224e-9 ua=-7.005982417e-10 lua=5.447513284e-16 ub=1.752388505e-18 lub=-1.139532890e-24 uc=3.570790382e-11 luc=2.928167858e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.603930204e+00 la0=-1.473840662e-6 ags=3.280924670e-01 lags=2.880340734e-7 a1=0.0 a2=0.42385546 b0=9.045966326e-08 lb0=8.103827942e-14 b1=5.181929613e-08 lb1=-3.422509015e-14 keta=5.571583279e-04 lketa=8.665127072e-9 dwg=0.0 dwb=0.0 pclm=1.111012835e+00 lpclm=-1.175322883e-6 pdiblc1=0.39 pdiblc2=2.515197032e-03 lpdiblc2=9.056794489e-9 pdiblcb=-3.713428750e-02 lpdiblcb=4.782712430e-8 drout=0.56 pscbe1=6.250038353e+08 lpscbe1=3.397526038e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593653295e-01 lkt1=-1.445527005e-7 kt2=-1.505275342e-02 lkt2=-6.448037594e-8 at=1.697338581e+05 lat=-1.171955854e-1 ute=-8.810097670e-01 lute=-1.649079246e-6 ua1=2.120317340e-09 lua1=-4.420641968e-15 pua1=-6.617444900e-36 ub1=-1.471838908e-18 lub1=3.150583117e-24 uc1=8.836977321e-12 luc1=9.269779387e-17 kt1l=0.0 prt=0.0 tvoff=3.291355927e-03 ltvoff=-4.669304753e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.148 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.337722202e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.210445684e-9 k1=5.909023591e-01 lk1=-3.456528306e-8 k2=-7.388526331e-02 lk2=3.200507309e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.776495273e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.902439363e-8 nfactor=3.165758097e+00 lnfactor=-8.184297285e-7 eta0=-1.412393438e-03 leta0=3.712885085e-09 weta0=1.734723476e-24 peta0=-1.734723476e-30 etab=7.846713825e-02 letab=-1.533135934e-07 wetab=-2.255140519e-23 petab=1.543903894e-28 u0=3.307948362e-02 lu0=-5.377884419e-9 ua=2.524868235e-10 lua=-1.305649982e-15 pua=1.654361225e-36 ub=3.598957487e-19 lub=1.563972301e-24 uc=6.136947818e-11 luc=-2.053990878e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.678388382e+04 lvsat=6.244044530e-3 a0=5.103841728e-01 la0=6.492636467e-7 ags=-2.518364953e-01 lags=1.413958035e-6 a1=0.0 a2=0.42385546 b0=2.064332386e-08 lb0=2.165857249e-13 b1=5.165556530e-08 lb1=-3.390720903e-14 keta=6.875730921e-02 lketa=-1.237445111e-07 wketa=-1.110223025e-22 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=1.622800558e-01 lpclm=6.666285246e-7 pdiblc1=4.235466902e-01 lpdiblc1=-6.513042940e-8 pdiblc2=9.520078457e-03 lpdiblc2=-4.543084728e-09 wpdiblc2=2.775557562e-23 pdiblcb=-2.408827873e-02 lpdiblcb=2.249848091e-8 drout=2.213441718e-01 ldrout=6.574955493e-7 pscbe1=8.622349078e+08 lpscbe1=-1.208282023e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.138758140e-06 lalpha0=1.003507157e-11 walpha0=1.270549421e-27 palpha0=5.188076802e-33 alpha1=0.85 beta0=1.046688446e+01 lbeta0=6.587686325e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.895211174e-01 lkt1=1.081429396e-7 kt2=-6.816647419e-02 lkt2=3.863916934e-8 at=1.533204212e+05 lat=-8.532912747e-2 ute=-2.347817386e+00 lute=1.198707212e-6 ua1=-1.510649725e-09 lua1=2.628829754e-15 pua1=8.271806126e-37 ub1=9.241642797e-19 lub1=-1.501223529e-24 pub1=7.703719778e-46 uc1=7.123910305e-11 luc1=-2.845505959e-17 kt1l=0.0 prt=0.0 tvoff=8.754564218e-04 ltvoff=2.113031463e-11 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.149 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.348772052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.170117734e-09 wvth0=-1.776356839e-21 k1=6.241244142e-01 lk1=-6.584338282e-8 k2=-6.309843653e-02 lk2=2.184942669e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.155802128e-01 ldsub=4.182060776e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.804439774e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.639345798e-8 nfactor=2.356259295e+00 lnfactor=-5.629793918e-8 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=3.747002708e-22 peta0=2.914335440e-28 etab=-1.583239050e-01 letab=6.962185877e-8 u0=3.145552919e-02 lu0=-3.848954058e-9 ua=-8.663853263e-10 lua=-2.522475177e-16 ub=1.918035997e-18 lub=9.700507105e-26 uc=2.808849155e-11 luc=1.079367420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.974950271e+04 lvsat=4.111139587e-2 a0=1.037003369e+00 la0=1.534590463e-7 ags=2.215750625e+00 lags=-9.092406929e-7 a1=0.0 a2=0.42385546 b0=4.720422507e-07 lb0=-2.084000451e-13 b1=2.945156505e-08 lb1=-1.300245365e-14 keta=-1.117400778e-01 lketa=4.619125183e-8 dwg=0.0 dwb=0.0 pclm=1.239890271e+00 lpclm=-3.479264066e-7 pdiblc1=6.380995512e-01 lpdiblc1=-2.671289443e-7 pdiblc2=8.798868557e-03 lpdiblc2=-3.864075704e-9 pdiblcb=8.317315894e-02 lpdiblcb=-7.848666099e-08 wpdiblcb=-7.632783294e-23 ppdiblcb=-7.199102425e-29 drout=8.488040648e-01 ldrout=6.675084452e-8 pscbe1=9.960958090e+08 lpscbe1=-2.468563667e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.950414640e-06 lalpha0=-1.346715358e-12 alpha1=0.85 beta0=1.697483351e+01 lbeta0=4.605434001e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.708668097e-01 lkt1=-3.568429924e-9 kt2=-1.865572788e-02 lkt2=-7.974505161e-9 at=1.086315090e+05 lat=-4.325514226e-02 pat=-1.164153218e-22 ute=-8.665203951e-01 lute=-1.959131673e-7 ua1=1.678807431e-09 lua1=-3.739995059e-16 ub1=-7.043401311e-19 lub1=3.199057490e-26 uc1=7.216247987e-11 luc1=-2.932440595e-17 kt1l=0.0 prt=0.0 tvoff=5.610461820e-04 ltvoff=3.171431537e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.150 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.234299035e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.292465884e-8 k1=1.440277361e-01 lk1=1.461125792e-7 k2=7.954110737e-02 lk2=-4.112393499e-08 wk2=-1.110223025e-22 pk2=-4.163336342e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.967001176e-01 ldsub=5.015590546e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-4.241165060e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.703595200e-8 nfactor=7.024742053e-01 lnfactor=6.738250248e-7 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.259628912e-02 letab=-1.466673405e-08 wetab=-1.040834086e-23 petab=-9.540979118e-30 u0=1.747213606e-02 lu0=2.324518243e-9 ua=-1.633387130e-09 lua=8.637304047e-17 ub=2.051759808e-18 lub=3.796788098e-26 uc=2.188162327e-11 luc=1.353391965e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.270649104e+05 lvsat=2.562865788e-3 a0=1.296210063e+00 la0=3.902291985e-8 ags=-6.815012499e-01 lags=3.698554483e-07 pags=3.330669074e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.112499912e-02 lketa=-2.571139951e-08 wketa=-5.551115123e-23 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=6.151398985e-01 lpclm=-7.210786358e-8 pdiblc1=-2.150883799e-01 lpdiblc1=1.095415826e-07 ppdiblc1=-2.775557562e-29 pdiblc2=-6.356604807e-03 lpdiblc2=2.826853609e-09 wpdiblc2=-4.770489559e-24 ppdiblc2=-1.301042607e-30 pdiblcb=-8.794872771e-02 lpdiblcb=-2.938743742e-9 drout=1.380423788e+00 ldrout=-1.679518208e-7 pscbe1=1.654406421e+08 lpscbe1=1.198662603e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.870637209e-06 lalpha0=-1.311494739e-12 alpha1=0.85 beta0=2.085046091e+01 lbeta0=-1.250491838e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-1.812142371e-01 lkt1=-4.314878560e-8 kt2=-4.272334130e-02 lkt2=2.651009219e-09 wkt2=1.110223025e-22 at=-3.181692230e+03 lat=6.108820692e-3 ute=-1.303565937e+00 lute=-2.963679176e-9 ua1=1.486947611e-09 lua1=-2.892960814e-16 ub1=-1.657962222e-18 lub1=4.530013775e-25 uc1=-1.025991505e-10 luc1=4.783040720e-17 wuc1=2.584939414e-32 puc1=1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=2.259348754e-03 ltvoff=-4.326336554e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.151 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.930860018e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.711422647e-8 k1=9.070734896e-01 lk1=4.493472261e-17 k2=-1.591041470e-01 lk2=4.573290196e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-6.810552122e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=4.755015826e-19 cit=0.0 voff='-1.280633099e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.654090323e-9 nfactor=5.957541296e+00 lnfactor=-3.324467521e-7 eta0=1.898829686e-03 leta0=-2.306811989e-10 etab=-4.399800002e-02 letab=1.940225758e-18 u0=2.922478324e-02 lu0=7.405084524e-11 ua=-1.220812587e-09 lua=7.370791619e-18 ub=2.115070575e-18 lub=2.584475532e-26 uc=1.195576603e-10 luc=-5.169673981e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.331606188e+05 lvsat=1.395622962e-3 a0=1.499999999e+00 la0=1.372715275e-16 ags=1.250000000e+00 lags=2.939160026e-17 a1=0.0 a2=0.42385546 b0=-6.354672333e-08 lb0=1.216830786e-14 b1=9.081564444e-11 lb1=-1.738992449e-17 keta=-1.805936561e-01 lketa=1.865947890e-08 pketa=-5.551115123e-29 dwg=0.0 dwb=0.0 pclm=3.411771752e-01 lpclm=-1.964783753e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.350031281e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301070776e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865729793e-18 drout=5.033266590e-01 ldrout=1.244684356e-16 pscbe1=7.914198799e+08 lpscbe1=1.229667664e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.021680590e-09 lalpha0=2.791544112e-15 alpha1=0.85 beta0=1.511289772e+01 lbeta0=-1.518288121e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.815303639e-01 lkt1=-4.791051739e-9 kt2=-2.887893901e-02 lkt2=7.457923168e-19 at=-1.466737011e+04 lat=8.308167207e-3 ute=-1.324741698e+00 lute=1.091182657e-9 ua1=-2.384733716e-11 lua1=1.407276948e-25 ub1=7.077531684e-19 lub1=1.999107579e-34 uc1=1.471862500e-10 luc1=-2.894304963e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.152 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-1.831149227e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.718331905e-08 wvth0=5.498473919e-07 pvth0=-6.679876025e-14 k1=0.90707349 k2=-3.177226182e-01 lk2=2.384321379e-08 wk2=7.808647454e-08 pk2=-9.486413446e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.116862511e+00 ldsub=-2.014520348e-07 wdsub=-9.461129123e-07 pdsub=1.149394733e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-7.534944890e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.870770867e-18 nfactor=1.481564214e+01 lnfactor=-1.408581992e-06 wnfactor=-5.815003466e-06 pnfactor=7.064415111e-13 eta0=-9.291641965e-03 leta0=1.128804440e-09 weta0=4.094194726e-09 peta0=-4.973873405e-16 etab=-0.043998 u0=1.023621911e-01 lu0=-8.811120290e-09 wu0=-3.770496766e-08 pu0=4.580625702e-15 ua=-2.719480416e-09 lua=1.894379515e-16 wua=7.047949674e-16 pua=-8.562272141e-23 ub=1.143211721e-17 lub=-1.106045972e-24 wub=-4.837085769e-24 pub=5.876382018e-31 uc=-1.483618842e-10 luc=2.737879980e-17 wuc=1.103154131e-16 puc=-1.340177828e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.397188281e+05 lvsat=5.988923570e-04 wvsat=1.109471491e-02 pvsat=-1.347852535e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-8.567887637e-06 lb0=1.045326668e-12 wb0=4.176588799e-12 pb0=-5.073970668e-19 b1=1.087199936e-08 lb1=-1.327152809e-15 wb1=-3.557169064e-14 pb1=4.321462409e-21 keta=-7.029957120e-01 lketa=8.212401507e-08 wketa=3.857447777e-07 pketa=-4.686259006e-14 dwg=0.0 dwb=0.0 pclm=2.588588800e-02 lpclm=1.865563978e-08 wpclm=1.156056326e-07 ppclm=-1.404446588e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000000e-08 lalpha0=-7.565063010e-26 walpha0=2.038405963e-22 palpha0=-2.476374937e-29 alpha1=0.85 beta0=1.390318600e+01 lbeta0=-4.865774312e-09 wbeta0=3.694822226e-17 pbeta0=-4.490630090e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=3.150525271e+00 lkt1=-4.338863625e-07 wkt1=-2.092985223e-06 pkt1=2.542684028e-13 kt2=-0.028878939 at=5.372048694e+04 lat=5.147885531e-12 wat=-2.407375723e-11 pat=2.924585715e-18 ute=-1.139353895e+00 lute=-2.143084008e-08 wute=-2.062934326e-07 pute=2.506176395e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.153 nmos lmin=2.0e-05 lmax=0.0001 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.154 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.708426337e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.252791506e-07 wvth0=1.261275650e-08 pvth0=-2.515171072e-13 k1=8.563148236e-01 lk1=-5.749272069e-06 wk1=-1.320090092e-07 pk1=2.632455809e-12 k2=-1.666668387e-01 lk2=2.443350368e-06 wk2=5.689881457e-08 pk2=-1.134646914e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.838467843e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.826312224e-07 wvoff=-2.057756625e-08 pvoff=4.103472492e-13 nfactor=2.665187130e+00 lnfactor=1.579821760e-06 wnfactor=4.686981286e-08 pnfactor=-9.346537170e-13 eta0=0.08 etab=-0.07 u0=2.114930307e-02 lu0=9.946208851e-08 wu0=1.798646804e-09 pu0=-3.586769007e-14 ua=-1.679070196e-09 lua=1.246374973e-14 wua=2.364472333e-16 pua=-4.715109193e-21 ub=2.294165355e-18 lub=-9.197718372e-24 wub=-1.847676444e-25 pub=3.684541394e-30 uc=6.319175009e-11 luc=-2.922374937e-16 wuc=2.680076753e-20 puc=-5.344471305e-25 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.005872261e+00 la0=7.113681217e-06 wa0=2.081000773e-07 pa0=-4.149824778e-12 ags=3.184325364e-01 lags=5.274017249e-07 wags=1.371568691e-09 pags=-2.735111785e-14 a1=0.0 a2=0.42385546 b0=1.544031141e-07 lb0=-1.640388914e-12 wb0=-4.538158201e-14 pb0=9.049761822e-19 b1=1.239155927e-07 lb1=-1.961556089e-12 wb1=-5.172232830e-14 pb1=1.031420086e-18 keta=-5.703606912e-03 lketa=2.307243714e-08 wketa=1.640837579e-09 pketa=-3.272073961e-14 dwg=0.0 dwb=0.0 pclm=6.813389444e-02 lpclm=-1.022178526e-06 wpclm=-4.202360349e-08 ppclm=8.380131006e-13 pdiblc1=0.39 pdiblc2=3.653257484e-03 lpdiblc2=-5.370102638e-08 wpdiblc2=-1.675864763e-09 ppdiblc2=3.341923372e-14 pdiblcb=-0.025 drout=0.56 pscbe1=-1.078769269e+08 lpscbe1=6.638060577e+03 wpscbe1=1.896089666e+01 ppscbe1=-3.781084552e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.038755871e-01 lkt1=3.488880050e-07 wkt1=1.116173142e-08 pkt1=-2.225815108e-13 kt2=-6.613201125e-02 lkt2=7.301391687e-07 wkt2=1.659377877e-08 pkt2=-3.309046070e-13 at=2.419035782e+05 lat=-1.334156769e+00 wat=-2.364773605e-02 pat=4.715709975e-7 ute=-5.424700958e-01 lute=-1.142507366e-05 wute=-2.561838073e-07 pute=5.108685806e-12 ua1=1.702128911e-09 lua1=-1.158857405e-14 wua1=-3.632292258e-16 pua1=7.243330521e-21 ub1=-9.722038958e-19 lub1=8.031112345e-24 wub1=3.182827621e-25 pub1=-6.347031245e-30 uc1=1.838810819e-10 luc1=-2.992473629e-15 wuc1=-6.202406092e-17 puc1=1.236851943e-21 kt1l=0.0 prt=0.0 tvoff=-9.125892064e-04 ltvoff=6.992859372e-08 wtvoff=1.404517870e-09 ptvoff=-2.800817344e-14 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.155 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.212948133e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=3.246138729e-07 wvth0=-4.370091234e-10 pvth0=-1.478825762e-13 k1=-3.097407272e-01 lk1=3.510941762e-06 wk1=4.039871954e-07 pk1=-1.624150546e-12 k2=3.252604521e-01 lk2=-1.463283325e-06 wk2=-1.705302161e-07 pk2=6.714775493e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.111747466e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.285420078e-07 wvoff=2.973757232e-08 pvoff=1.077028075e-14 nfactor=2.582618861e+00 lnfactor=2.235536508e-06 wnfactor=1.833238696e-07 pnfactor=-2.018301698e-12 eta0=0.08 etab=-0.07 u0=3.314519519e-02 lu0=4.196879213e-09 wu0=-3.170652976e-09 pu0=3.595934570e-15 ua=1.446953856e-10 lua=-2.019659107e-15 wua=-6.056346203e-16 pua=1.972272058e-21 ub=8.090157013e-19 lub=2.596576810e-24 wub=5.567113138e-25 pub=-2.203903372e-30 uc=-9.056390868e-11 luc=9.288109178e-16 wuc=5.423022578e-17 puc=-4.309901880e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.302931750e+00 la0=-3.186898555e-06 wa0=-4.834592548e-07 pa0=1.342183977e-12 ags=1.619529349e-01 lags=1.770082289e-06 wags=1.076895562e-07 pags=-8.716739270e-13 a1=0.0 a2=0.42385546 b0=-3.627311905e-07 lb0=2.466425926e-12 wb0=2.171236131e-13 pb0=-1.179705150e-18 b1=-1.763186854e-07 lb1=4.227502265e-13 wb1=9.539642161e-14 pb1=-1.369214070e-19 keta=-9.571346744e-03 lketa=5.378803887e-08 wketa=-4.219481527e-09 pketa=1.381890252e-14 dwg=0.0 dwb=0.0 pclm=-2.214557099e+00 lpclm=1.710578004e-05 wpclm=8.252993143e-07 ppclm=-6.049819708e-12 pdiblc1=0.39 pdiblc2=-4.258106338e-03 lpdiblc2=9.126958658e-09 wpdiblc2=1.428780577e-09 ppdiblc2=8.763736215e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.130084801e+09 lpscbe1=-3.193195151e+03 wpscbe1=-2.653204113e+02 ppscbe1=1.879507572e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.014860218e-01 lkt1=3.299113056e-07 wkt1=8.203734939e-09 pkt1=-1.990906232e-13 kt2=2.884516595e-02 lkt2=-2.412075437e-08 wkt2=-2.094096326e-08 pkt2=-3.282297866e-14 at=8.777267782e+03 lat=5.172125619e-01 wat=7.094320816e-02 pat=-2.796216618e-7 ute=-3.090541061e+00 lute=8.810396234e-06 wute=1.005164263e-06 pute=-4.908292236e-12 ua1=-2.326505799e-09 lua1=2.040477210e-14 wua1=2.076114407e-15 pua1=-1.212868279e-20 ub1=1.868921578e-18 lub1=-1.453164583e-23 wub1=-1.565041819e-24 pub1=8.609364552e-30 uc1=-3.308670284e-10 luc1=1.095391283e-15 wuc1=1.406259684e-16 puc1=-3.724904283e-22 kt1l=0.0 prt=0.0 tvoff=1.170616184e-02 ltvoff=-3.028304106e-08 wtvoff=-3.192691262e-09 ptvoff=8.500498518e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.156 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.754813741e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.110383021e-07 wvth0=-2.484661161e-08 pvth0=-5.167246974e-14 k1=7.204051047e-01 lk1=-5.493636122e-07 wk1=-8.711361213e-08 pk1=3.115164118e-13 k2=-8.321597051e-02 lk2=1.467207760e-07 wk2=2.578014226e-08 pk2=-1.022769800e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.134444189e+00 ldsub=-6.205649728e-06 wdsub=-6.937504918e-07 pdsub=2.734407851e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.101285257e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.244183425e-07 wvoff=3.323818981e-08 pvoff=-3.027354079e-15 nfactor=1.958702583e+00 lnfactor=4.694693785e-06 wnfactor=2.089383660e-07 pnfactor=-2.119260877e-12 eta0=4.972277100e-01 leta0=-1.644497178e-06 weta0=-1.838438803e-07 peta0=7.246180805e-13 etab=-4.347462371e-01 letab=1.437642187e-06 wetab=1.607188639e-07 petab=-6.334711521e-13 u0=3.417493305e-02 lu0=1.381818520e-10 wu0=-2.384585909e-09 pu0=4.976622288e-16 ua=-1.618969024e-09 lua=4.931799471e-15 wua=4.965006326e-16 pua=-2.371778611e-21 ub=3.422017333e-18 lub=-7.702532541e-24 wub=-9.026547728e-25 pub=3.548167627e-30 uc=2.138032809e-10 luc=-2.708480989e-16 wuc=-9.628405992e-17 puc=1.622597619e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.708634921e+05 lvsat=-1.146434382e+00 wvsat=-1.572501115e-01 pvsat=6.197991128e-7 a0=4.927508956e+00 la0=-1.353163287e-05 wa0=-1.796833028e-06 pa0=6.518828316e-12 ags=-1.483012567e-01 lags=2.992944842e-06 wags=2.575536916e-07 pags=-1.462361319e-12 a1=0.0 a2=0.42385546 b0=2.131173423e-07 lb0=1.967269960e-13 wb0=-6.631266636e-14 pb0=-6.254502224e-20 b1=-1.289456209e-07 lb1=2.360299561e-13 wb1=9.772729862e-14 pb1=-1.461085262e-19 keta=5.835703204e-02 lketa=-2.139507151e-07 wketa=-3.124846132e-08 pketa=1.203532480e-13 dwg=0.0 dwb=0.0 pclm=9.223100401e+00 lpclm=-2.797558687e-05 wpclm=-4.385654125e-06 ppclm=1.448908032e-11 pdiblc1=0.39 pdiblc2=1.587233328e-02 lpdiblc2=-7.021688725e-08 wpdiblc2=-7.221295281e-09 ppdiblc2=4.285788911e-14 pdiblcb=-9.060184120e-02 lpdiblcb=2.585687387e-07 wpdiblcb=2.890627049e-08 ppdiblcb=-1.139336604e-13 drout=0.56 pscbe1=-1.460852652e+08 lpscbe1=1.836811297e+03 wpscbe1=4.168754426e+02 ppscbe1=-8.093578355e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-5.462624123e-02 lkt1=-6.430830634e-07 wkt1=-1.106885027e-07 pkt1=2.695214672e-13 kt2=1.678743451e-01 lkt2=-5.721023175e-07 wkt2=-9.889624312e-08 pkt2=2.744366655e-13 at=3.007507517e+05 lat=-6.335968372e-01 wat=-7.083192521e-02 pat=2.791830416e-7 ute=2.328061426e+00 lute=-1.254694961e-05 wute=-1.734926577e-06 pute=5.891737449e-12 ua1=1.282642596e-08 lua1=-3.932029627e-14 wua1=-5.788064913e-15 pua1=1.886786991e-20 ub1=-8.190206301e-18 lub1=2.511626588e-23 wub1=3.632164400e-24 pub1=-1.187535100e-29 uc1=-2.078670485e-10 luc1=6.105885843e-16 wuc1=1.171571309e-16 puc1=-2.799883338e-22 kt1l=0.0 prt=0.0 tvoff=7.093315405e-03 ltvoff=-1.210157141e-08 wtvoff=-2.055460956e-09 ptvoff=4.018121190e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.157 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.433558434e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.073902984e-08 wvth0=-5.924441339e-08 pvth0=1.511038085e-14 k1=4.579373377e-01 lk1=-3.978611713e-08 wk1=7.188514544e-08 pk1=2.822549961e-15 k2=-7.831836337e-02 lk2=1.372121403e-07 wk2=2.396675750e-09 pk2=-5.687830719e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-2.306442577e+00 ldsub=2.416269756e-06 wdsub=1.387500984e-06 pdsub=-1.306312751e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.181522212e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.415236497e-08 wvoff=2.189705241e-08 pvoff=1.899130541e-14 nfactor=6.055486354e+00 lnfactor=-3.259154551e-06 wnfactor=-1.562279567e-06 pnfactor=1.319533942e-12 eta0=-6.815196765e-01 leta0=6.440243706e-07 weta0=3.676877606e-07 peta0=-3.461728790e-13 etab=1.021758658e+00 letab=-1.390141675e-06 wetab=-5.099735807e-07 petab=6.686688394e-13 u0=3.208826625e-02 lu0=4.189416225e-09 wu0=5.358838294e-10 pu0=-5.172388881e-15 ua=2.480366747e-09 lua=-3.027003537e-15 wua=-1.204463179e-15 pua=9.306188149e-22 ub=-3.331521713e-18 lub=5.409368968e-24 wub=1.995698405e-24 pub=-2.078944491e-30 uc=1.194050659e-10 luc=-8.757528605e-17 wuc=-3.137589587e-17 puc=3.624147009e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.208594326e+05 lvsat=-1.917612078e-01 wvsat=1.068523015e-01 pvsat=1.070479756e-7 a0=-3.850179839e+00 la0=3.510127038e-06 wa0=2.357460443e-06 pa0=-1.546674297e-12 ags=-2.818333424e+00 lags=8.176774914e-06 wags=1.387530367e-06 pags=-3.656195215e-12 a1=0.0 a2=0.42385546 b0=-1.163262504e-06 lb0=2.868949199e-12 wb0=6.400573758e-13 pb0=-1.433952570e-18 b1=-3.010178232e-09 lb1=-8.471942723e-15 wb1=2.955405026e-14 pb1=-1.375111889e-20 keta=2.921957431e-01 lketa=-6.679452989e-07 wketa=-1.207979674e-07 pketa=2.942123604e-13 dwg=0.0 dwb=0.0 pclm=-1.020372996e+01 lpclm=9.741332307e-06 wpclm=5.604196729e-06 ppclm=-4.906075255e-12 pdiblc1=1.398595626e+00 lpdiblc1=-1.958174287e-06 wpdiblc1=-5.271426560e-07 ppdiblc1=1.023440087e-12 pdiblc2=-3.907636767e-02 lpdiblc2=3.646524634e-08 wpdiblc2=2.627279386e-08 ppdiblc2=-2.217041604e-14 pdiblcb=-2.007094305e-02 lpdiblcb=1.216339873e-07 wpdiblcb=-2.171900223e-09 ppdiblcb=-5.359582710e-14 drout=-8.799957498e-01 ldrout=2.795731588e-06 wdrout=5.954196045e-07 pdrout=-1.155998826e-12 pscbe1=1.136461827e+09 lpscbe1=-6.532359265e+02 wpscbe1=-1.482558477e+02 ppscbe1=2.878366528e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.791396051e-05 lalpha0=5.425280811e-11 walpha0=1.231300321e-11 palpha0=-2.390552334e-17 alpha1=0.85 beta0=-4.484268428e+00 lbeta0=3.561514033e-05 wbeta0=8.083071686e-06 pbeta0=-1.569317052e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-5.789964456e-01 lkt1=3.749743472e-07 wkt1=1.024364257e-07 pkt1=-1.442575976e-13 kt2=-2.178706246e-01 lkt2=1.768161408e-07 wkt2=8.093485427e-08 pkt2=-7.470289242e-14 at=1.705295737e+05 lat=-3.807742432e-01 wat=-9.303818512e-03 pat=1.597270838e-7 ute=-5.540609384e+00 lute=2.729964609e-06 wute=1.726125523e-06 pute=-8.278467493e-13 ua1=-1.183785219e-08 lua1=8.565054442e-15 wua1=5.583216121e-15 pua1=-3.209313025e-21 ub1=6.973487581e-18 lub1=-4.323833504e-24 wub1=-3.270457755e-24 pub1=1.525993276e-30 uc1=1.955596937e-10 luc1=-1.726587877e-16 wuc1=-6.721168955e-17 puc1=7.796114994e-23 kt1l=0.0 prt=0.0 tvoff=-5.404607971e-04 ltvoff=2.719298209e-09 wtvoff=7.654901579e-10 ptvoff=-1.458715905e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.158 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.011662335e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.898189724e-08 wvth0=-3.583796993e-08 pvth0=-6.926457976e-15 k1=7.543784998e-01 lk1=-3.188813210e-07 wk1=-7.041952680e-08 pk1=1.368004066e-13 k2=-1.480453023e-02 lk2=7.741475564e-08 wk2=-2.610923115e-08 pk2=-3.004039492e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.958005786e-01 ldsub=6.044285648e-08 wdsub=1.069350322e-08 pdsub=-1.006778357e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.525610920e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.175689477e-08 wvoff=3.898881994e-08 pvoff=2.899645558e-15 nfactor=3.325124673e+00 lnfactor=-6.885572539e-07 wnfactor=-5.237996271e-07 pnfactor=3.418196179e-13 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=-1.734723476e-23 peta0=5.117434254e-29 etab=-8.545727191e-01 letab=3.763980475e-07 wetab=3.764143889e-07 petab=-1.658530245e-13 u0=5.826424875e-02 lu0=-2.045490483e-08 wu0=-1.449365167e-08 pu0=8.977708379e-15 ua=9.430879384e-10 lua=-1.579677061e-15 wua=-9.782591500e-16 pua=7.176508887e-22 ub=1.673851876e-18 lub=6.968798093e-25 wub=1.320137499e-25 pub=-3.243114795e-31 uc=-1.839725578e-10 luc=1.980504994e-16 wuc=1.146469892e-16 puc=-1.012370319e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.423027942e+05 lvsat=1.108732169e-01 wvsat=2.606128974e-01 pvsat=-3.771547285e-8 a0=-1.003107947e+00 la0=8.296487113e-07 wa0=1.102949461e-06 pa0=-3.655697710e-13 ags=1.037681674e+01 lags=-4.246274235e-06 wags=-4.412133497e-06 pags=1.804107118e-12 a1=0.0 a2=0.42385546 b0=4.900328083e-06 lb0=-2.839836449e-12 wb0=-2.394073026e-12 pb0=1.422638726e-18 b1=-1.439010381e-09 lb1=-9.951175258e-15 wb1=1.670043358e-14 pb1=-1.649618739e-21 keta=-7.585476610e-01 lketa=3.213149057e-07 wketa=3.496848773e-07 pketa=-1.487406512e-13 dwg=0.0 dwb=0.0 pclm=5.292984057e-01 lpclm=-3.636636405e-07 wpclm=3.841687014e-07 ppclm=8.508052220e-15 pdiblc1=5.035810452e-01 lpdiblc1=-1.115530590e-06 wpdiblc1=7.272500894e-08 ppdiblc1=4.586730783e-13 pdiblc2=4.284342353e-03 lpdiblc2=-4.358255090e-09 wpdiblc2=2.440697331e-09 ppdiblc2=2.671691894e-16 pdiblcb=5.598187126e-01 lpdiblcb=-4.243240050e-07 wpdiblcb=-2.576898390e-07 ppdiblcb=1.869707350e-13 drout=3.051484297e+00 ldrout=-9.057018350e-07 wdrout=-1.190839419e-06 pdrout=5.257390370e-13 pscbe1=1.860156694e+09 lpscbe1=-1.334584512e+03 wpscbe1=-4.671389645e+02 ppscbe1=5.880606428e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.966165067e-05 lalpha0=-9.368683756e-12 walpha0=-1.768474096e-11 palpha0=4.336932819e-18 alpha1=0.85 beta0=3.746953021e+01 lbeta0=-3.883773732e-06 wbeta0=-1.108008887e-05 pbeta0=2.348676860e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-1.985287990e-01 lkt1=1.676938451e-08 wkt1=-3.910824340e-08 pkt1=-1.099527329e-14 kt2=-7.540427180e-02 lkt2=4.268606410e-08 wkt2=3.068007880e-08 pkt2=-2.738872488e-14 at=-4.913103341e+05 lat=2.423387642e-01 wat=3.243477585e-01 pat=-1.544012048e-7 ute=-4.493789002e+00 lute=1.744397875e-06 wute=1.961017482e-06 pute=-1.048994239e-12 ua1=-7.657055565e-09 lua1=4.628892954e-15 wua1=5.047266283e-15 pua1=-2.704723756e-21 ub1=7.705763646e-18 lub1=-5.013261167e-24 wub1=-4.546771225e-24 pub1=2.727624540e-30 uc1=4.091688214e-10 luc1=-3.737687909e-16 wuc1=-1.821964124e-16 puc1=1.862176567e-22 kt1l=0.0 prt=0.0 tvoff=2.350099521e-03 ltvoff=-2.123862560e-12 wtvoff=-9.672194849e-10 ptvoff=1.726059655e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.159 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='7.917397333e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.515363489e-08 wvth0=-9.099367987e-08 pvth0=1.742401578e-14 k1=-6.381025958e-01 lk1=2.958795879e-07 wk1=4.228446856e-07 pk1=-8.096883746e-14 k2=3.870867572e-01 lk2=-1.000146213e-07 wk2=-1.662690198e-07 pk2=3.183818952e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.362593861e-01 ldsub=4.258085937e-08 wdsub=-2.138700644e-08 pdsub=4.095312315e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380513e-03 lcdscd=-1.132138095e-9 cit=0.0 voff='-5.729250391e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.553070277e-08 wvoff=8.045065487e-08 pvoff=-1.540517410e-14 nfactor=-1.156010523e-01 lnfactor=8.304749836e-07 wnfactor=4.422776627e-07 pnfactor=-8.468998052e-14 eta0=8.647808876e-01 leta0=-1.654605149e-7 etab=3.016462838e-02 letab=-1.420110506e-08 wetab=1.314633609e-09 petab=-2.517339312e-16 u0=-1.608969592e-03 lu0=5.978282839e-09 wu0=1.031585631e-08 pu0=-1.975342061e-15 ua=-3.747676847e-09 lua=4.912299213e-16 wua=1.143052678e-15 pua=-2.188785852e-22 ub=4.020043276e-18 lub=-3.389308473e-25 wub=-1.064117028e-24 pub=2.037635133e-31 uc=3.964209863e-10 luc=-5.818512481e-17 wuc=-2.024879649e-16 puc=3.877361045e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.451651668e+05 lvsat=1.121369143e-01 wvsat=3.093658911e-01 pvsat=-5.923923702e-8 a0=3.982463849e-01 la0=2.109703927e-07 wa0=4.854678991e-07 pa0=-9.296030612e-14 ags=3.823503236e-01 lags=1.661427659e-07 wags=-5.751522039e-07 pags=1.101335949e-13 a1=0.0 a2=0.42385546 b0=-2.705640818e-06 lb0=5.180923377e-13 wb0=1.462756007e-12 pb0=-2.800972967e-19 b1=-4.234591278e-08 lb1=8.108649455e-15 wb1=2.289355552e-14 pb1=-4.383795372e-21 keta=9.393643650e-03 lketa=-1.772042917e-08 wketa=2.256130617e-08 pketa=-4.320174273e-15 dwg=0.0 dwb=0.0 pclm=-7.026744782e-01 lpclm=1.802351402e-07 wpclm=7.124526221e-07 ppclm=-1.364247028e-13 pdiblc1=-3.846247109e+00 lpdiblc1=8.048576431e-07 wpdiblc1=1.963120606e-06 ppdiblc1=-3.759101124e-13 pdiblc2=-1.630572281e-02 lpdiblc2=4.731970419e-09 wpdiblc2=5.378811564e-09 ppdiblc2=-1.029967111e-15 pdiblcb=-6.295687482e-01 lpdiblcb=1.007739075e-07 wpdiblcb=2.928171149e-07 ppdiblcb=-5.607037807e-14 drout=1.380423010e+00 ldrout=-1.679516718e-07 wdrout=4.206827544e-13 pdrout=-8.055485790e-20 pscbe1=-2.659588805e+09 lpscbe1=6.608198490e+02 wpscbe1=1.527301320e+03 ppscbe1=-2.924568205e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.254897462e-05 lalpha0=-6.228536856e-12 walpha0=-1.388253091e-11 palpha0=2.658310314e-18 alpha1=0.85 beta0=3.966567905e+01 lbeta0=-4.853342698e-06 wbeta0=-1.017210901e-05 pbeta0=1.947816466e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=2.788189658e-02 lkt1=-8.318776785e-08 wkt1=-1.130440609e-07 pkt1=2.164635505e-14 kt2=5.970418509e-02 lkt2=-1.696242810e-08 wkt2=-5.537559845e-08 pkt2=1.060365184e-14 at=7.973023548e+04 lat=-9.767652698e-03 wat=-4.482484130e-02 pat=8.583329562e-9 ute=5.212499897e-02 lute=-2.625595137e-07 wute=-7.329299021e-07 pute=1.403458152e-13 ua1=5.011906208e-09 lua1=-9.642763031e-16 wua1=-1.905705416e-15 pua1=3.649159072e-22 ub1=-6.987196886e-18 lub1=1.473475206e-24 wub1=2.881154795e-24 pub1=-5.517008071e-31 uc1=-8.852423636e-10 luc1=1.976956255e-16 wuc1=4.231219656e-16 puc1=-8.102193270e-23 kt1l=0.0 prt=0.0 tvoff=4.141648699e-03 ltvoff=-7.930677427e-10 wtvoff=-1.017631584e-09 ptvoff=1.948622015e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.160 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='3.188721406e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.539388895e-08 wvth0=1.482487882e-07 pvth0=-2.838756746e-14 k1=9.070734896e-01 lk1=4.493605488e-17 k2=-1.235937631e-01 lk2=-2.226451182e-09 wk2=-1.919804989e-08 pk2=3.676157781e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.721187889e+00 ldsub=-2.417621599e-07 wdsub=-6.825791966e-07 pdsub=1.307043600e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=7.733163068e-19 wcdscd=8.408412855e-19 pcdscd=-1.610092268e-25 cit=0.0 voff='-5.788064174e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.665690436e-08 wvoff=2.436861477e-07 pvoff=-4.666248568e-14 nfactor=6.034329297e+00 lnfactor=-3.471505793e-07 wnfactor=-4.151405086e-08 pnfactor=7.949359543e-15 eta0=1.898828344e-03 leta0=-2.306809055e-10 weta0=8.284599205e-16 peta0=-1.586384763e-22 etab=-4.399800002e-02 letab=1.940225758e-18 u0=-2.157061589e-02 lu0=9.800658642e-09 wu0=2.746161822e-08 pu0=-5.258515426e-15 ua=-1.216624623e-09 lua=6.568855202e-18 wua=-2.264147192e-18 pua=4.335524892e-25 ub=3.059510342e-18 lub=-1.550022378e-25 wub=-5.105943599e-25 pub=9.777167161e-32 uc=2.300983891e-10 luc=-2.633667597e-17 wuc=-5.976185527e-17 puc=1.144355862e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.907304479e+05 lvsat=-4.792539333e-02 wvsat=-1.392504918e-01 pvsat=2.666451968e-8 a0=1.499999999e+00 la0=1.372710834e-16 ags=1.250000000e+00 lags=2.939071209e-17 a1=0.0 a2=0.42385546 b0=7.842042470e-06 lb0=-1.501641344e-12 wb0=-4.274014497e-12 pb0=8.184139399e-19 b1=1.257296856e-07 lb1=-2.407547457e-14 wb1=-6.792439352e-14 pb1=1.300657042e-20 keta=-4.970054985e-01 lketa=7.924791697e-08 wketa=1.710623672e-07 pketa=-3.275604845e-14 dwg=0.0 dwb=0.0 pclm=3.541932009e-01 lpclm=-2.214022424e-08 wpclm=-7.036880037e-09 ppclm=1.347464011e-15 pdiblc1=3.569721502e-01 lpdiblc1=-2.350042383e-17 pdiblc2=8.406112095e-03 lpdiblc2=6.301018735e-19 pdiblcb=-1.032957700e-01 lpdiblcb=1.865702037e-18 drout=5.033266590e-01 ldrout=1.244683245e-16 pscbe1=7.914198799e+08 lpscbe1=1.229643822e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.722018768e-07 lalpha0=-2.883815094e-14 walpha0=-8.930169984e-14 palpha0=1.710002530e-20 alpha1=0.85 beta0=1.921843729e+01 lbeta0=-9.379821624e-07 wbeta0=-2.219586069e-06 pbeta0=4.250196581e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=1.147967078e+00 lkt1=-2.976683989e-07 wkt1=-8.268952611e-07 pkt1=1.583388660e-13 kt2=-2.887893901e-02 lkt2=7.458408890e-19 at=-9.113968307e+04 lat=2.295154453e-02 wat=4.134337950e-02 pat=-7.916678367e-9 ute=-1.043961853e+00 lute=-5.267422672e-08 wute=-1.517985691e-07 pute=2.906730080e-14 ua1=-2.384733716e-11 lua1=1.407276883e-25 ub1=7.077531684e-19 lub1=1.999107579e-34 uc1=1.471862500e-10 luc1=-2.894563457e-27 kt1l=0.0 prt=0.0 tvoff=1.179891318e-02 ltvoff=-2.259326690e-09 wtvoff=-6.378870033e-09 ptvoff=1.221464307e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.161 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='1.684958986e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.405665375e-07 wvth0=-4.600931415e-07 pvth0=4.551746021e-14 k1=0.90707349 k2=-5.992990256e-02 lk2=-9.960718943e-09 wk2=-6.128451691e-08 pk2=8.789074314e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-7.650469660e-01 ldsub=6.028056767e-08 wdsub=6.119395721e-07 pdsub=-2.656154709e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000004e-03 lcdscd=-4.073512361e-19 wcdscd=-1.961961843e-18 pcdscd=1.794920549e-25 cit=0.0 voff='-1.029050771e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.884155414e-08 wvoff=-5.656358136e-08 pvoff=-1.018634709e-14 nfactor=3.673279571e+00 lnfactor=-6.031609237e-08 wnfactor=2.089142965e-07 pnfactor=-2.247417866e-14 eta0=-9.291641602e-03 leta0=1.128804616e-09 weta0=4.094195032e-09 peta0=-4.973874356e-16 etab=-0.043998 u0=1.113089050e-01 lu0=-6.342342828e-09 wu0=-4.254184746e-08 pu0=3.245925605e-15 ua=-2.636320704e-09 lua=1.790420532e-16 wua=6.598361659e-16 pua=-8.000236614e-23 ub=8.689859253e-18 lub=-8.390108056e-25 wub=-3.354533364e-24 pub=4.432704455e-31 uc=-4.137594320e-10 luc=5.188303529e-17 wuc=2.537978202e-16 puc=-2.664955212e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.913281879e+05 lvsat=7.138098211e-02 wvsat=4.063221253e-01 pvsat=-3.961491528e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-2.701428726e-05 lb0=2.732914729e-12 wb0=1.414930272e-11 pb0=-1.419761176e-18 b1=-2.822838249e-07 lb1=2.549245476e-14 wb1=1.229177289e-13 pb1=-1.017807567e-20 keta=3.529876863e-02 lketa=1.458040076e-08 wketa=-1.340084400e-08 pketa=-1.034635077e-14 dwg=0.0 dwb=0.0 pclm=-4.484420980e-03 lpclm=2.143408533e-08 wpclm=1.320247935e-07 ppclm=-1.554658246e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.554204558e-07 lalpha0=3.526057576e-14 walpha0=2.083706321e-13 palpha0=-1.906299562e-20 alpha1=0.85 beta0=4.323593680e+00 lbeta0=8.715328080e-07 wbeta0=5.179034154e-06 pbeta0=-4.738091184e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.192225113e+00 lkt1=2.296041896e-07 wkt1=1.336108602e-06 pkt1=-1.044358214e-13 kt2=-0.028878939 at=2.321558836e+05 lat=-1.632434069e-02 wat=-9.646788540e-02 pat=8.825460961e-9 ute=-1.780539257e+00 lute=3.680961573e-08 wute=1.403518923e-07 pute=-6.424890150e-15 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-1.512313749e-02 ltvoff=1.011325558e-09 wtvoff=8.176052066e-09 ptvoff=-5.467549590e-16 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.162 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.163 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.994668746e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.544692521e-7 k1=5.567246685e-01 lk1=2.250008142e-7 k2=-3.753682867e-02 lk2=-1.316939191e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.305469020e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.863852027e-8 nfactor=2.771556646e+00 lnfactor=-5.413444673e-07 wnfactor=-3.552713679e-21 eta0=0.08 etab=-0.07 u0=2.523127352e-02 lu0=1.806153189e-8 ua=-1.142460886e-09 lua=1.762962689e-15 ub=1.874841192e-18 lub=-8.357714558e-25 uc=6.325257356e-11 luc=-2.934504041e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.478148621e+00 la0=-2.304211214e-6 ags=3.215452670e-01 lags=4.653292520e-7 a1=0.0 a2=0.42385546 b0=5.141108901e-08 lb0=4.134251128e-13 b1=6.533449983e-09 lb1=3.792182659e-13 keta=-1.979779367e-03 lketa=-5.118621772e-8 dwg=0.0 dwb=0.0 pclm=-2.723730757e-02 lpclm=8.796649638e-7 pdiblc1=0.39 pdiblc2=-1.500631174e-04 lpdiblc2=2.214283815e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.484578828e+07 lpscbe1=5.779955729e+03 ppscbe1=3.814697266e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.785444005e-01 lkt1=-1.562534981e-7 kt2=-2.847296976e-02 lkt2=-2.083808001e-8 at=1.882358100e+05 lat=-2.639417198e-1 ute=-1.123870918e+00 lute=1.689227007e-7 ua1=8.777919913e-10 lua1=4.849929102e-15 ub1=-2.498715138e-19 lub1=-6.373268737e-24 uc1=4.311949195e-11 luc1=-1.854783527e-16 kt1l=0.0 prt=0.0 tvoff=2.274918442e-03 ltvoff=6.364954573e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.164 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.203030353e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.100082638e-8 k1=6.070950799e-01 lk1=-1.750151033e-7 k2=-6.175232989e-02 lk2=6.061314481e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.436862930e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.529848099e-7 nfactor=2.998666424e+00 lnfactor=-2.344933585e-6 eta0=0.08 etab=-0.07 u0=2.594950133e-02 lu0=1.235773582e-8 ua=-1.229772697e-09 lua=2.456348214e-15 ub=2.072453931e-18 lub=-2.405110249e-24 uc=3.250982582e-11 luc=-4.930730334e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.205736687e+00 la0=-1.408556515e-7 ags=4.063508819e-01 lags=-2.081533517e-7 a1=0.0 a2=0.42385546 b0=1.300237912e-07 lb0=-2.108765609e-13 b1=4.018039235e-08 lb1=1.120115442e-13 keta=-1.914732290e-02 lketa=8.514958892e-08 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=-3.415671334e-01 lpclm=3.375910875e-06 ppclm=-1.332267630e-27 pdiblc1=0.39 pdiblc2=-1.015535266e-03 lpdiblc2=2.901597311e-08 ppdiblc2=1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=5.279487523e+08 lpscbe1=1.072286184e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.828679120e-01 lkt1=-1.219183917e-7 kt2=-1.867966943e-02 lkt2=-9.861143742e-8 at=1.697805725e+05 lat=-1.173797096e-1 ute=-8.093534416e-01 lute=-2.328813438e-6 ua1=2.385168358e-09 lua1=-7.120879208e-15 ub1=-1.682889954e-18 lub1=5.007027145e-24 uc1=-1.172096455e-11 luc1=2.500363649e-16 kt1l=0.0 prt=0.0 tvoff=4.460452809e-03 ltvoff=-1.099143601e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.165 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.190927967e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.230688184e-9 k1=5.227035938e-01 lk1=1.576127577e-7 k2=-2.470877571e-02 lk2=-8.539350536e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.346955344e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.175478609e-7 nfactor=2.432881412e+00 lnfactor=-1.148998834e-7 eta0=0.08 etab=-0.07 u0=2.876319284e-02 lu0=1.267610102e-9 ua=-4.921769782e-10 lua=-4.508749862e-16 ub=1.373471670e-18 lub=3.499185461e-25 uc=-4.710263065e-12 luc=9.739515593e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.398947600e+04 lvsat=2.601795562e-1 a0=8.496548100e-01 la0=1.262636082e-6 ags=4.362084739e-01 lags=-3.258366324e-7 a1=0.0 a2=0.42385546 b0=6.262290173e-08 lb0=5.478310126e-14 b1=9.284330643e-08 lb1=-9.555859435e-14 keta=-1.256033512e-02 lketa=5.918706878e-08 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=-7.299990678e-01 lpclm=4.906909907e-6 pdiblc1=0.39 pdiblc2=-5.161616168e-04 lpdiblc2=2.704769886e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.058302000e-01 lkt1=-3.141285524e-8 kt2=-5.656746377e-02 lkt2=5.072277354e-8 at=140000.0 ute=-1.609298042e+00 lute=8.241570060e-7 ua1=-3.093992072e-10 lua1=3.499721124e-15 ub1=5.287273135e-20 lub1=-1.834457180e-24 uc1=5.801725153e-11 luc1=-2.483583746e-17 kt1l=0.0 prt=0.0 tvoff=2.428513583e-03 ltvoff=-2.982575995e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.166 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.089025731e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.355348830e-8 k1=6.210783384e-01 lk1=-3.338043174e-8 k2=-7.287918567e-02 lk2=8.128671184e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.684575726e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.105221472e-8 nfactor=2.509943663e+00 lnfactor=-2.645151643e-7 eta0=1.529357436e-01 leta0=-1.416037250e-7 etab=-1.356098056e-01 letab=1.273805191e-7 u0=3.330443718e-02 lu0=-7.549152198e-9 ua=-2.531232828e-10 lua=-9.149943890e-16 ub=1.197650942e-18 lub=6.912720282e-25 uc=4.819849020e-11 luc=-5.326447822e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.216383920e+05 lvsat=5.118069287e-2 a0=1.5 ags=3.306216395e-01 lags=-1.208412716e-7 a1=0.0 a2=0.42385546 b0=2.893269030e-07 lb0=-3.853595433e-13 b1=6.406177809e-08 lb1=-3.967966003e-14 keta=1.804868298e-02 lketa=-2.399113257e-10 dwg=0.0 dwb=0.0 pclm=2.514812332e+00 lpclm=-1.392845999e-6 pdiblc1=2.022625040e-01 lpdiblc1=3.644897201e-7 pdiblc2=2.054888393e-02 lpdiblc2=-1.384979216e-8 pdiblcb=-0.025 drout=4.712896868e-01 ldrout=1.722298312e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.465203076e-01 lkt1=4.758641904e-8 kt2=-3.419160390e-02 lkt2=7.280354855e-9 at=1.494148600e+05 lat=-1.827881888e-2 ute=-1.623223622e+00 lute=8.511933232e-7 ua1=8.330753023e-10 lua1=1.281622859e-15 ub1=-4.487099786e-19 lub1=-8.606413705e-25 uc1=4.302494914e-11 luc1=4.271507725e-18 kt1l=0.0 prt=0.0 tvoff=1.196794232e-03 ltvoff=-5.912101179e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.167 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.198331257e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.262526024e-9 k1=5.945636729e-01 lk1=-8.417245317e-9 k2=-7.405858157e-02 lk2=9.239055919e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.200691365e-01 ldsub=3.759434895e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.640772326e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.517624344e-8 nfactor=2.136378447e+00 lnfactor=8.719125697e-8 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=1.387778781e-22 peta0=5.724587471e-29 etab=-0.0003125 u0=2.537137744e-02 lu0=-8.028751188e-11 ua=-1.277039402e-09 lua=4.900830196e-17 ub=1.973452790e-18 lub=-3.913455073e-26 uc=7.621505733e-11 luc=-3.170365354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.491497045e+05 lvsat=2.527917735e-2 a0=1.5 ags=3.636231996e-01 lags=-1.519117784e-7 a1=0.0 a2=0.42385546 b0=-5.329428236e-07 lb0=3.887958925e-13 b1=3.646208073e-08 lb1=-1.369493136e-14 keta=3.505080060e-02 lketa=-1.624716703e-8 dwg=0.0 dwb=0.0 pclm=1.401156785e+00 lpclm=-3.443548925e-7 pdiblc1=6.686280889e-01 lpdiblc1=-7.458694891e-8 pdiblc2=9.823425603e-03 lpdiblc2=-3.751923299e-9 pdiblcb=-0.025 drout=3.489129465e-01 ldrout=2.874458189e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.732940400e-07 lalpha0=4.738442925e-13 walpha0=-1.588186776e-28 palpha0=-2.646977960e-35 alpha1=0.85 beta0=1.232362872e+01 lbeta0=1.446472051e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.872836861e-01 lkt1=-8.184030794e-9 kt2=-5.776830313e-03 lkt2=-1.947175667e-8 at=2.447863600e+05 lat=-1.080697509e-1 ute=-4.332357624e-02 lute=-6.362604508e-7 ua1=3.797551190e-09 lua1=-1.509389686e-15 ub1=-2.612985844e-18 lub1=1.176994057e-24 uc1=-4.320013795e-12 luc1=4.884612750e-17 kt1l=0.0 prt=0.0 tvoff=1.550263425e-04 ltvoff=3.895997652e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.168 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-6.460861841e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.179995785e-07 wvth0=5.425584298e-07 pvth0=-2.395319509e-13 k1=3.215296738e-01 lk1=1.121234428e-07 wk1=-6.246443363e-16 pk1=2.757716278e-22 k2=2.027032227e-01 lk2=-1.129474060e-07 wk2=-8.502373418e-08 pk2=3.753678831e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.918636815e+00 ldsub=-7.122995012e-07 wdsub=-7.626963377e-07 pdsub=3.367197554e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380526e-03 lcdscd=-1.132138101e-09 wcdscd=-5.670290626e-18 pcdscd=2.503351693e-24 cit=0.0 voff='-1.312856297e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.478450304e-07 wvoff=4.064880447e-07 pvoff=-1.794587809e-13 nfactor=-9.494418017e+00 lnfactor=5.222025065e-06 wnfactor=4.574884540e-06 pnfactor=-2.019747476e-12 eta0=8.575034974e-01 leta0=-1.622476491e-07 weta0=3.206650982e-09 peta0=-1.415691515e-15 etab=3.314814668e-02 letab=-1.477240706e-08 wetab=-2.697061064e-17 petab=1.190713598e-23 u0=-4.549974592e-02 lu0=3.120832125e-08 wu0=2.965553687e-08 pu0=-1.309250435e-14 ua=-9.152852427e-10 lua=-1.107010946e-16 wua=-1.049896989e-16 pua=4.635148220e-23 ub=3.715186442e-18 lub=-8.080855737e-25 wub=-9.297873515e-25 pub=4.104880987e-31 uc=-7.466179277e-11 luc=3.490636351e-17 wuc=5.086182201e-18 puc=-2.245478235e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.540764798e+05 lvsat=-1.976389250e-01 wvsat=-1.749951541e-01 pvsat=7.725791062e-8 a0=1.500000005e+00 la0=-2.051548265e-15 wa0=-1.908173175e-15 pa0=8.424314579e-22 ags=-9.229389053e-01 lags=4.160873790e-07 wags=-4.085576322e-16 pags=1.803725294e-22 a1=0.0 a2=0.42385546 b0=1.183614983e-05 lb0=-5.071985346e-12 wb0=-4.944822290e-12 pb0=2.183069813e-18 b1=1.813073448e-07 lb1=-7.764208762e-14 wb1=-7.565522668e-14 pb1=3.340072341e-20 keta=2.154659923e-01 lketa=-9.589794835e-08 wketa=-6.824076496e-08 pketa=3.012734236e-14 dwg=0.0 dwb=0.0 pclm=3.122201696e-01 lpclm=1.363953781e-07 wpclm=2.652575637e-07 ppclm=-1.171075007e-13 pdiblc1=6.089912889e-01 lpdiblc1=-4.825813664e-08 wpdiblc1=3.266755755e-16 ppdiblc1=-1.442224118e-22 pdiblc2=-4.098684799e-03 lpdiblc2=2.394493534e-09 wpdiblc2=-8.758905060e-18 ppdiblc2=3.866935418e-24 pdiblcb=3.497017532e-02 lpdiblcb=-2.647599282e-08 wpdiblcb=-2.593453230e-17 ppdiblcb=1.144969536e-23 drout=1.380423969e+00 ldrout=-1.679518564e-07 wdrout=-1.730208865e-15 pdrout=7.638623067e-22 pscbe1=8.065718918e+08 lpscbe1=-2.901398245e+00 wpscbe1=-1.709299088e-07 ppscbe1=7.546329498e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.357543124e-06 lalpha0=-3.344446835e-13 walpha0=-1.385880676e-13 palpha0=6.118469163e-20 alpha1=0.85 beta0=1.741913130e+01 lbeta0=-8.031210008e-07 wbeta0=-3.695681838e-07 pbeta0=1.631591792e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=1.717064543e+00 lkt1=-8.930757130e-07 wkt1=-8.573519888e-07 pkt1=3.785089001e-13 kt2=-6.596893542e-02 lkt2=7.102215049e-09 wkt2=-1.036781772e-17 pkt2=4.577241364e-24 at=1.352622736e+05 lat=-5.971640012e-02 wat=-6.929403432e-02 pat=3.059234604e-8 ute=-1.191874099e+00 lute=-1.291914746e-07 wute=-1.847840914e-07 pute=8.157958940e-14 ua1=6.869697213e-10 lua1=-1.361115162e-16 wua1=-1.956225900e-24 pua1=8.636461461e-31 ub1=-4.485097332e-19 lub1=2.214081566e-25 wub1=-2.778912954e-33 pub1=1.226850994e-39 uc1=7.501918240e-11 luc1=1.381898313e-17 wuc1=4.023675333e-26 puc1=-1.776396215e-32 kt1l=0.0 prt=0.0 tvoff=1.800798793e-02 ltvoff=-7.492232833e-09 wtvoff=-7.127584371e-09 ptvoff=3.146728714e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.169 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.052884800e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.732735793e-07 wvth0=-1.937708678e-06 pvth0=2.354044764e-13 k1=9.070734846e-01 lk1=6.600062719e-16 wk1=2.230873264e-15 pk1=-2.710198732e-22 k2=-8.563009731e-01 lk2=8.983707145e-08 wk2=3.036561935e-07 pk2=-3.688997632e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-6.009741069e+00 ldsub=8.058738663e-07 wdsub=2.723915492e-06 pdsub=-3.309175974e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999951e-03 lcdscd=5.991289062e-18 wcdscd=2.025101614e-17 pcdscd=-2.460215191e-24 cit=0.0 voff='3.268914957e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.295000199e-07 wvoff=-1.451743017e-06 pvoff=1.763664522e-13 nfactor=4.302065645e+01 lnfactor=-4.833876484e-06 wnfactor=-1.633887336e-05 pnfactor=1.984944369e-12 eta0=2.788951197e-02 leta0=-3.388184913e-09 weta0=-1.145232494e-08 peta0=1.391297147e-15 etab=-4.399800023e-02 letab=2.849745440e-17 wetab=9.632361575e-17 petab=-1.170195885e-23 u0=2.811179085e-01 lu0=-3.133438692e-08 wu0=-1.059126317e-07 pu0=1.286690197e-14 ua=-2.072729848e-09 lua=1.109333431e-16 wua=3.749632103e-16 pua=-4.555278056e-23 ub=-5.635417563e-18 lub=9.824241847e-25 wub=3.320669113e-24 pub=-4.034148078e-31 uc=1.356955340e-10 luc=-5.374119570e-18 wuc=-1.816493643e-17 puc=2.206785467e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.343671922e+06 lvsat=1.849019255e-01 wvsat=6.249826933e-01 pvsat=-7.592664748e-8 a0=1.499999983e+00 la0=2.016197875e-15 wa0=6.814900644e-15 pa0=-8.279155139e-22 ags=1.249999996e+00 lags=4.316866864e-16 wags=1.459135035e-15 pags=-1.772644254e-22 a1=0.0 a2=0.42385546 b0=-4.193667106e-05 lb0=5.224757035e-12 wb0=1.766007961e-11 pb0=-2.145452431e-18 b1=-6.416263659e-07 lb1=7.993819691e-14 wb1=2.701972381e-13 pb1=-3.282518167e-20 keta=-6.618928660e-01 lketa=7.210398998e-08 wketa=2.437170177e-07 pketa=-2.960820561e-14 dwg=0.0 dwb=0.0 pclm=2.488199722e+00 lpclm=-2.802742426e-07 wpclm=-9.473484416e-07 ppclm=1.150895728e-13 pdiblc1=3.569721528e-01 lpdiblc1=-3.451687824e-16 wpdiblc1=-1.166696961e-15 ppdiblc1=1.417373996e-22 pdiblc2=8.406112024e-03 lpdiblc2=9.254763622e-18 wpdiblc2=3.128181048e-17 ppdiblc2=-3.800300352e-24 pdiblcb=-1.032957702e-01 lpdiblcb=2.740263572e-17 wpdiblcb=9.262302036e-17 ppdiblcb=-1.125241567e-23 drout=5.033266450e-01 ldrout=1.828157625e-15 wdrout=6.179313061e-15 pdrout=-7.506999467e-22 pscbe1=7.914198785e+08 lpscbe1=1.806063652e-07 wpscbe1=6.104640961e-07 ppscbe1=-7.416296005e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.153755122e-06 lalpha0=1.464337724e-13 walpha0=4.949573845e-13 palpha0=-6.013039281e-20 alpha1=0.85 beta0=1.118571965e+01 lbeta0=3.904900632e-07 wbeta0=1.319886371e-06 pbeta0=-1.603477156e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-7.677689364e+00 lkt1=9.058881336e-07 wkt1=3.061971388e-06 pkt1=-3.719866561e-13 kt2=-2.887893909e-02 lkt2=1.095470936e-17 wkt2=3.702776974e-17 pkt2=-4.498360018e-24 at=-5.589570783e+05 lat=7.321688670e-02 wat=2.474786940e-01 pat=-3.006519662e-8 ute=-2.886183374e+00 lute=1.952450311e-07 wute=6.599431837e-07 pute=-8.017385762e-14 ua1=-2.384735301e-11 lua1=2.066970792e-24 wua1=6.986519862e-24 pua1=-8.487643461e-31 ub1=7.077531458e-19 lub1=2.936231578e-33 wub1=9.924688323e-33 pub1=-1.205710723e-39 uc1=1.471862503e-10 luc1=-4.251460194e-26 wuc1=-1.437023655e-25 puc1=1.745785362e-32 kt1l=0.0 prt=0.0 tvoff=-6.044851437e-02 ltvoff=7.531088967e-09 wtvoff=2.545565847e-08 ptvoff=-3.092506125e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.170 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-3.435598678e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.579583245e-07 wvth0=1.796188423e-06 pvth0=-2.182117468e-13 k1=0.90707349 k2=-2.107921637e+00 lk2=2.418914594e-07 wk2=8.411261769e-07 pk2=-1.021850547e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.948957557e+00 ldsub=-2.824825950e-07 wdsub=-1.024569669e-06 pdsub=1.244708708e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='2.710812388e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.616983712e-07 wvoff=-1.296377536e-06 pvoff=1.574917213e-13 nfactor=-9.718055751e+00 lnfactor=1.573138706e-06 wnfactor=6.109565162e-06 pnfactor=-7.422266333e-13 eta0=4.841478680e-04 leta0=-5.881718202e-11 weta0=-2.133310221e-10 peta0=2.591673255e-17 etab=-0.043998 u0=2.649207452e-01 lu0=-2.936665834e-08 wu0=-1.102281398e-07 pu0=1.339117580e-14 ua=-3.027207701e-09 lua=2.268890396e-16 wua=8.320734854e-16 pua=-1.010852794e-22 ub=1.372746819e-17 lub=-1.369895353e-24 wub=-5.574265064e-24 pub=6.771951656e-31 uc=-1.088917355e-10 luc=2.433980945e-17 wuc=1.194633573e-16 puc=-1.451312543e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.613456549e+05 lvsat=-8.297683985e-02 wvsat=-2.337724555e-01 pvsat=2.840008053e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-4.381579665e-06 lb0=6.623392016e-13 wb0=4.176607507e-12 pb0=-5.073993396e-19 b1=7.740561823e-08 lb1=-7.414122714e-15 wb1=-3.557294977e-14 pb1=4.321615375e-21 keta=-8.705490917e-01 lketa=9.745280022e-08 wketa=3.857447104e-07 pketa=-4.686258189e-14 dwg=0.0 dwb=0.0 pclm=3.277891720e-02 lpclm=1.802500936e-08 wpclm=1.156053743e-07 ppclm=-1.404443450e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.174699132e-07 lalpha0=-8.002272280e-15 walpha0=2.976834824e-21 palpha0=-3.616437609e-28 alpha1=0.85 beta0=1.607724329e+01 lbeta0=-2.037615779e-07 wbeta0=2.059408644e-14 pbeta0=-2.501892027e-21 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.409528512e+00 lkt1=2.658803443e-07 wkt1=9.912274339e-07 pkt1=-1.204202560e-13 kt2=-0.028878939 at=1.322515441e+04 lat=3.704755975e-03 wat=-3.293820191e-10 pat=4.001532216e-17 ute=-9.550152712e-01 lute=-3.936485696e-08 wute=-2.234003926e-07 pute=2.714002010e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=-3.511084150e-02 ltvoff=4.452916439e-09 wtvoff=1.698327406e-08 ptvoff=-2.063230032e-15 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.171 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.507213+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.044140846 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.32810784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.74441 eta0=0.08 etab=-0.07 u0=0.026137 ua=-1.0540541e-9 ub=1.83293e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=7.2143e-8 b1=2.555e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0025941 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.172 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='4.994668746e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.544692521e-7 k1=5.567246685e-01 lk1=2.250008142e-7 k2=-3.753682867e-02 lk2=-1.316939191e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.305469020e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.863852027e-8 nfactor=2.771556646e+00 lnfactor=-5.413444673e-7 eta0=0.08 etab=-0.07 u0=2.523127352e-02 lu0=1.806153189e-08 wu0=-2.775557562e-23 ua=-1.142460886e-09 lua=1.762962689e-15 ub=1.874841192e-18 lub=-8.357714558e-25 uc=6.325257356e-11 luc=-2.934504041e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.478148621e+00 la0=-2.304211214e-6 ags=3.215452670e-01 lags=4.653292520e-7 a1=0.0 a2=0.42385546 b0=5.141108901e-08 lb0=4.134251128e-13 b1=6.533449983e-09 lb1=3.792182659e-13 keta=-1.979779367e-03 lketa=-5.118621772e-8 dwg=0.0 dwb=0.0 pclm=-2.723730757e-02 lpclm=8.796649638e-07 ppclm=2.220446049e-28 pdiblc1=0.39 pdiblc2=-1.500631174e-04 lpdiblc2=2.214283815e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.484578828e+07 lpscbe1=5.779955729e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.785444005e-01 lkt1=-1.562534981e-7 kt2=-2.847296976e-02 lkt2=-2.083808001e-8 at=1.882358100e+05 lat=-2.639417198e-1 ute=-1.123870918e+00 lute=1.689227007e-7 ua1=8.777919913e-10 lua1=4.849929102e-15 ub1=-2.498715138e-19 lub1=-6.373268737e-24 uc1=4.311949195e-11 luc1=-1.854783527e-16 kt1l=0.0 prt=0.0 tvoff=2.274918442e-03 ltvoff=6.364954573e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.173 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.203030353e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.100082638e-8 k1=6.070950799e-01 lk1=-1.750151033e-7 k2=-6.175232989e-02 lk2=6.061314481e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.436862930e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.529848099e-7 nfactor=2.998666424e+00 lnfactor=-2.344933585e-6 eta0=0.08 etab=-0.07 u0=2.594950133e-02 lu0=1.235773582e-8 ua=-1.229772697e-09 lua=2.456348214e-15 ub=2.072453931e-18 lub=-2.405110249e-24 uc=3.250982582e-11 luc=-4.930730334e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.205736687e+00 la0=-1.408556515e-7 ags=4.063508819e-01 lags=-2.081533517e-07 wags=-4.440892099e-22 a1=0.0 a2=0.42385546 b0=1.300237912e-07 lb0=-2.108765609e-13 b1=4.018039235e-08 lb1=1.120115442e-13 keta=-1.914732290e-02 lketa=8.514958892e-8 dwg=0.0 dwb=0.0 pclm=-3.415671334e-01 lpclm=3.375910875e-06 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.015535266e-03 lpdiblc2=2.901597311e-08 ppdiblc2=-1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=5.279487523e+08 lpscbe1=1.072286184e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.828679120e-01 lkt1=-1.219183917e-7 kt2=-1.867966943e-02 lkt2=-9.861143742e-8 at=1.697805725e+05 lat=-1.173797096e-1 ute=-8.093534416e-01 lute=-2.328813438e-6 ua1=2.385168358e-09 lua1=-7.120879208e-15 ub1=-1.682889954e-18 lub1=5.007027145e-24 uc1=-1.172096455e-11 luc1=2.500363649e-16 kt1l=0.0 prt=0.0 tvoff=4.460452809e-03 ltvoff=-1.099143601e-8 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.174 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.190927967e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.230688184e-9 k1=5.227035938e-01 lk1=1.576127577e-7 k2=-2.470877571e-02 lk2=-8.539350536e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.346955344e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.175478609e-7 nfactor=2.432881412e+00 lnfactor=-1.148998834e-7 eta0=0.08 etab=-0.07 u0=2.876319284e-02 lu0=1.267610102e-9 ua=-4.921769782e-10 lua=-4.508749862e-16 ub=1.373471670e-18 lub=3.499185461e-25 uc=-4.710263065e-12 luc=9.739515593e-17 puc=5.169878828e-38 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.398947600e+04 lvsat=2.601795562e-1 a0=8.496548100e-01 la0=1.262636082e-6 ags=4.362084739e-01 lags=-3.258366324e-7 a1=0.0 a2=0.42385546 b0=6.262290173e-08 lb0=5.478310126e-14 b1=9.284330642e-08 lb1=-9.555859435e-14 keta=-1.256033512e-02 lketa=5.918706878e-08 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=-7.299990678e-01 lpclm=4.906909907e-06 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=-5.161616168e-04 lpdiblc2=2.704769886e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.058302000e-01 lkt1=-3.141285524e-8 kt2=-5.656746377e-02 lkt2=5.072277354e-08 wkt2=5.551115123e-23 at=140000.0 ute=-1.609298042e+00 lute=8.241570060e-07 wute=1.776356839e-21 ua1=-3.093992072e-10 lua1=3.499721124e-15 ub1=5.287273135e-20 lub1=-1.834457180e-24 uc1=5.801725153e-11 luc1=-2.483583746e-17 kt1l=0.0 prt=0.0 tvoff=2.428513583e-03 ltvoff=-2.982575995e-9 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.175 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.089025731e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.355348830e-8 k1=6.210783384e-01 lk1=-3.338043174e-8 k2=-7.287918567e-02 lk2=8.128671184e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.424458000e-01 ldsub=-5.483645665e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.684575726e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.105221472e-8 nfactor=2.509943663e+00 lnfactor=-2.645151643e-7 eta0=1.529357436e-01 leta0=-1.416037250e-7 etab=-1.356098056e-01 letab=1.273805191e-7 u0=3.330443718e-02 lu0=-7.549152198e-9 ua=-2.531232828e-10 lua=-9.149943890e-16 ub=1.197650942e-18 lub=6.912720282e-25 uc=4.819849020e-11 luc=-5.326447822e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.216383920e+05 lvsat=5.118069287e-2 a0=1.5 ags=3.306216395e-01 lags=-1.208412716e-7 a1=0.0 a2=0.42385546 b0=2.893269030e-07 lb0=-3.853595433e-13 pb0=2.117582368e-34 b1=6.406177809e-08 lb1=-3.967966003e-14 keta=1.804868298e-02 lketa=-2.399113257e-10 dwg=0.0 dwb=0.0 pclm=2.514812332e+00 lpclm=-1.392845999e-6 pdiblc1=2.022625040e-01 lpdiblc1=3.644897201e-7 pdiblc2=2.054888393e-02 lpdiblc2=-1.384979216e-8 pdiblcb=-0.025 drout=4.712896868e-01 ldrout=1.722298312e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.465203076e-01 lkt1=4.758641904e-8 kt2=-3.419160390e-02 lkt2=7.280354855e-9 at=1.494148600e+05 lat=-1.827881888e-2 ute=-1.623223622e+00 lute=8.511933232e-7 ua1=8.330753023e-10 lua1=1.281622859e-15 ub1=-4.487099786e-19 lub1=-8.606413705e-25 uc1=4.302494914e-11 luc1=4.271507725e-18 kt1l=0.0 prt=0.0 tvoff=1.196794232e-03 ltvoff=-5.912101179e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.176 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='5.198331257e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.262526024e-9 k1=5.945636729e-01 lk1=-8.417245317e-9 k2=-7.405858157e-02 lk2=9.239055919e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.200691365e-01 ldsub=3.759434895e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.640772326e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.517624344e-8 nfactor=2.136378447e+00 lnfactor=8.719125697e-8 eta0=-4.278900071e-01 leta0=4.052355877e-07 weta0=-1.110223025e-22 peta0=-1.474514955e-28 etab=-0.0003125 u0=2.537137744e-02 lu0=-8.028751188e-11 ua=-1.277039402e-09 lua=4.900830196e-17 ub=1.973452790e-18 lub=-3.913455073e-26 uc=7.621505733e-11 luc=-3.170365354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.491497045e+05 lvsat=2.527917735e-2 a0=1.5 ags=3.636231996e-01 lags=-1.519117784e-7 a1=0.0 a2=0.42385546 b0=-5.329428236e-07 lb0=3.887958925e-13 pb0=2.117582368e-34 b1=3.646208073e-08 lb1=-1.369493136e-14 wb1=-2.646977960e-29 keta=3.505080060e-02 lketa=-1.624716703e-8 dwg=0.0 dwb=0.0 pclm=1.401156785e+00 lpclm=-3.443548925e-7 pdiblc1=6.686280889e-01 lpdiblc1=-7.458694891e-8 pdiblc2=9.823425603e-03 lpdiblc2=-3.751923299e-9 pdiblcb=-0.025 drout=3.489129465e-01 ldrout=2.874458189e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.732940400e-07 lalpha0=4.738442925e-13 walpha0=1.058791184e-28 palpha0=-2.646977960e-35 alpha1=0.85 beta0=1.232362872e+01 lbeta0=1.446472051e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-2.872836861e-01 lkt1=-8.184030794e-9 kt2=-5.776830313e-03 lkt2=-1.947175667e-8 at=2.447863600e+05 lat=-1.080697509e-1 ute=-4.332357624e-02 lute=-6.362604508e-7 ua1=3.797551190e-09 lua1=-1.509389686e-15 ub1=-2.612985844e-18 lub1=1.176994057e-24 uc1=-4.320013795e-12 luc1=4.884612750e-17 puc1=-2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=1.550263425e-04 ltvoff=3.895997652e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.177 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='6.751903598e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.532551779e-8 k1=3.215296722e-01 lk1=1.121234435e-7 k2=-4.352569801e-03 lk2=-2.153517240e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=6.126491588e-02 ldsub=1.077041891e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.964380512e-03 lcdscd=-1.132138095e-09 wcdscd=6.938893904e-24 cit=0.0 voff='-3.229479487e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.081435351e-8 nfactor=1.646663388e+00 lnfactor=3.033935994e-7 eta0=8.653125600e-01 leta0=-1.656952409e-7 etab=3.314814661e-02 letab=-1.477240703e-08 wetab=1.301042607e-23 petab=-3.252606517e-31 u0=2.671950846e-02 lu0=-6.754684848e-10 ua=-1.170963560e-09 lua=2.177303096e-18 ub=1.450902724e-18 lub=1.915639877e-25 uc=-6.227556325e-11 luc=2.943801658e-17 wuc=-6.462348536e-33 puc=8.077935669e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.279159416e+05 lvsat=-9.495013609e-03 wvsat=2.328306437e-16 a0=1.5 ags=-9.229389063e-01 lags=4.160873794e-07 wags=3.885780586e-22 pags=-1.873501354e-28 a1=0.0 a2=0.42385546 b0=-2.058300694e-07 lb0=2.443801911e-13 pb0=1.058791184e-34 b1=-2.933597640e-09 lb1=3.697709100e-15 pb1=-1.654361225e-36 keta=4.928126982e-02 lketa=-2.252971997e-08 wketa=2.081668171e-23 pketa=3.469446952e-30 dwg=0.0 dwb=0.0 pclm=9.581940919e-01 lpclm=-1.487930650e-7 pdiblc1=6.089912897e-01 lpdiblc1=-4.825813699e-8 pdiblc2=-4.098684820e-03 lpdiblc2=2.394493543e-09 ppdiblc2=-4.336808690e-31 pdiblcb=3.497017526e-02 lpdiblcb=-2.647599279e-8 drout=1.380423965e+00 ldrout=-1.679518545e-7 pscbe1=8.065718914e+08 lpscbe1=-2.901398061e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.020043690e-06 lalpha0=-1.854434083e-13 alpha1=0.85 beta0=1.651913280e+01 lbeta0=-4.057842633e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-3.708194719e-01 lkt1=2.869584913e-8 kt2=-6.596893545e-02 lkt2=7.102215060e-9 at=-3.348744469e+04 lat=1.478423801e-2 ute=-1.641873348e+00 lute=6.947689369e-8 ua1=6.869697165e-10 lua1=-1.361115141e-16 ub1=-4.485097400e-19 lub1=2.214081596e-25 wub1=9.629649722e-41 pub1=2.407412430e-47 uc1=7.501918250e-11 luc1=1.381898309e-17 kt1l=0.0 prt=0.0 tvoff=6.503919024e-04 ltvoff=1.709028056e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.178 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='0.33404+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.90707349 k2=-0.116816 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.62373 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.266472+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.23108 eta0=0.0 etab=-0.043998 u0=0.023192 ua=-1.159593e-9 ub=2.45131e-18 uc=9.1459e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=178330.0 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=1.0704e-6 b1=1.6377e-8 keta=-0.068376 dwg=0.0 dwb=0.0 pclm=0.18115 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.16e-8 alpha1=0.85 beta0=14.4 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=43720.487 ute=-1.2790432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0015429 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.179 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-1.0316e-8 lint=2.9257e-8 vth0='-3.531268488e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.348115179e-08 wvth0=5.304268509e-07 pvth0=-6.443943641e-14 k1=0.90707349 k2=-4.094792879e-01 lk2=3.555449219e-08 wk2=1.436913983e-07 pk2=-1.745649321e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.018083006e+00 ldsub=-2.908803693e-07 wdsub=-1.052954790e-06 pdsub=1.279192657e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-4.462175937e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.183657320e-8 nfactor=-2.972044984e+00 lnfactor=7.535928418e-07 wnfactor=3.339437269e-06 pnfactor=-4.056948761e-13 eta0=7.747629855e-04 leta0=-9.412284665e-11 weta0=-3.326668770e-10 peta0=4.041436822e-17 etab=-0.043998 u0=6.530240354e-02 lu0=-5.115824484e-09 wu0=-2.825846097e-08 pu0=3.433007390e-15 ua=-2.717298978e-09 lua=1.892394685e-16 wua=7.048150466e-16 pua=-8.562516075e-23 ub=1.193222840e-17 lub=-1.151798852e-24 wub=-4.837082158e-24 pub=5.876377631e-31 uc=-1.169516676e-10 luc=2.531897836e-17 wuc=1.227730234e-16 puc=-1.491520352e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.513622016e+05 lvsat=-8.872390042e-03 wvsat=1.670626994e-02 pvsat=-2.029577910e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=-4.381559583e-06 lb0=6.623367619e-13 wb0=4.176599261e-12 pb0=-5.073983378e-19 b1=7.740263310e-08 lb1=-7.413760063e-15 wb1=-3.557172398e-14 pb1=4.321466459e-21 keta=-8.705488195e-01 lketa=9.745276715e-08 wketa=3.857445986e-07 pketa=-4.686256831e-14 dwg=0.0 dwb=0.0 pclm=3.277875141e-02 lpclm=1.802502951e-08 wpclm=1.156054423e-07 ppclm=-1.404444277e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.174699199e-07 lalpha0=-8.002273094e-15 walpha0=2.268604107e-22 palpha0=-2.756037423e-29 alpha1=0.85 beta0=1.607724334e+01 lbeta0=-2.037615840e-07 wbeta0=3.967670636e-17 pbeta0=-4.824585176e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=2.3267e-8 dwc=-3.2175e-8 xpart=0.0 cgso=2.4083264e-10 cgdo=2.4083264e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001041645846 mjs=0.44 pbsws=0.2 cjsws=2.856175336e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=1.852257592e-10 mjswgs=0.8 tnom=30.0 kt1=3.391387185e-01 lkt1=-6.804424281e-08 wkt1=-1.374632882e-07 pkt1=1.669986504e-14 kt2=-0.028878939 at=1.322515368e+04 lat=3.704756064e-03 wat=-2.678728197e-11 pat=3.254273906e-18 ute=-9.399429465e-01 lute=-4.119593340e-08 wute=-2.295895715e-07 pute=2.789191868e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=6.248024980e-03 ltvoff=-5.716068133e-10 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.ends sky130_fd_pr__nfet_01v8