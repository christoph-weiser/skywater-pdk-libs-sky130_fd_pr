* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.model sky130_fd_pr__diode_pd2nw_05v5_hvt d level=3.0 tlevc=1.0 area=1.0e+12 cj='0.00075561*1e-12*sky130_fd_pr__pfet_01v8_hvt__ajunction_mult' mj=0.34629 pb=0.6587 cjsw='9.2435e-011*1e-6*sky130_fd_pr__pfet_01v8_hvt__pjunction_mult' mjsw=0.26859 php=0.7418 cta=0.0012407 ctp=0 tpb=0.0019551 tphp=0.00014242 js=2.17e-017 jsw=8.2e-016 n=1.2556 rs=600 ik='4.76e-008/1e-12' ikr='0/1e-12' vb=12.8 ibv=0.00106 trs=0 eg=1.05 xti=2.0 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0