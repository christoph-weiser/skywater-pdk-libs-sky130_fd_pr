* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_top c0 c1 m5 sub
xsky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_0[0|0] c0 c1 m5 sub sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
xsky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_0[1|0] c0 c1 m5 sub sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
xsky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_0[0|1] c0 c1 m5 sub sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
xsky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5_0[1|1] c0 c1 m5 sub sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5
.ends