* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_03v3_nvt__toxe_mult=1.052
.param sky130_fd_pr__nfet_03v3_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__overlap_mult=1.37
.param sky130_fd_pr__nfet_03v3_nvt__ajunction_mult=1.3878
.param sky130_fd_pr__nfet_03v3_nvt__pjunction_mult=1.2464
.param sky130_fd_pr__nfet_03v3_nvt__lint_diff=-1.7325e-8
.param sky130_fd_pr__nfet_03v3_nvt__wint_diff=3.2175e-8
.param sky130_fd_pr__nfet_03v3_nvt__dlc_diff=-3.0000e-8
.param sky130_fd_pr__nfet_03v3_nvt__dwc_diff=3.2175e-8
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_0=0.070007
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_0=0.025405
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0=-1.8
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0=0.01866
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_0=-0.0034806
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0=-4720.5
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_0=-1.0e-18
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_0=1.1794e-11
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_1=7.2867e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_1=0.061113
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_1=0.022045
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1=-1.5295
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1=0.030601
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_1=-0.00236
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1=937.82
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_1=-7.7567e-19
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_2=4.3331e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_2=8.8389e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_2=0.0117
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2=-0.4369
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2=0.057242
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_2=0.011419
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2=5633.8
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_3=-2.5164e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_3=9.4843e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_3=0.077321
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_3=0.024946
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3=-1.8358
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3=0.012417
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_3=-0.0043072
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3=-3550.1
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_4=4.2773e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_4=1.029e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_4=0.017434
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_4=0.0092175
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4=-1.2004
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4=0.076144
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_4=0.0014096
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4=-4990.9
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_5=0.0070104
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5=-3975.1
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_5=4.2056e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_5=1.6413e-10
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_5=0.021544
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5=-1.6491
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5=0.10543
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6=-0.70119
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6=0.059414
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_6=0.0049892
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6=2172.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_6=2.8836e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_6=2.4441e-10
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_6=0.020119
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_7=0.069322
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_7=0.021677
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7=-1.4753
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7=0.028831
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_7=-0.0053542
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7=-1407.8
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_7=-4.6026e-19
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_7=-2.6093e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_8=0.013898
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8=-0.33169
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8=0.050109
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_8=0.0080728
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8=4767.8
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_8=3.6297e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_8=-2.7576e-13
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8=0.0
.include "sky130_fd_pr__nfet_03v3_nvt.pm3.spice"