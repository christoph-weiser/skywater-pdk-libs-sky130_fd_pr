* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_pfet_01v8__toxe_slope=1.267e-02
.param sky130_fd_pr__rf_pfet_01v8__toxe1_slope=1.067e-02
.param sky130_fd_pr__rf_pfet_01v8__toxe2_slope=1.167e-02
.param sky130_fd_pr__rf_pfet_01v8__toxe3_slope=1.367e-02
.param sky130_fd_pr__rf_pfet_01v8__toxe4_slope=1.467e-02
.param sky130_fd_pr__rf_pfet_01v8__toxe5_slope=1.567e-02
.param sky130_fd_pr__rf_pfet_01v8__nfactor_slope=0.429
.param sky130_fd_pr__rf_pfet_01v8__nfactor1_slope=0.0
.param sky130_fd_pr__rf_pfet_01v8__b_toxe_slope=6.443e-03
.param sky130_fd_pr__rf_pfet_01v8__b_toxe_slope1=4.443e-03
.param sky130_fd_pr__rf_pfet_01v8__b_nfactor_slope1=0.1
.param sky130_fd_pr__rf_pfet_01v8__b_voff_slope=0.014
.param sky130_fd_pr__rf_pfet_01v8__b_voff_slope1=0.009
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope1=7.356e-03
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope2=9.356e-03
.param sky130_fd_pr__rf_pfet_01v8__b_vth0_slope3=8.356e-03