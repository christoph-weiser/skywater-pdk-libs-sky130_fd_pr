* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_lvt__toxe_mult=1.052
.param sky130_fd_pr__pfet_01v8_lvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_lvt__overlap_mult=0.10000
.param sky130_fd_pr__pfet_01v8_lvt__ajunction_mult=1.0909e+0
.param sky130_fd_pr__pfet_01v8_lvt__pjunction_mult=1.0909e+0
.param sky130_fd_pr__pfet_01v8_lvt__lint_diff=-1.7325e-8
.param sky130_fd_pr__pfet_01v8_lvt__wint_diff=3.2175e-8
.param sky130_fd_pr__pfet_01v8_lvt__dlc_diff=-5.9781e-8
.param sky130_fd_pr__pfet_01v8_lvt__dwc_diff=3.2175e-8
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_0=0.00013132
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_0=0.42229
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0=-0.17989
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_0=-0.080656
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_0=-0.050109
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_1=-0.03983
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_1=4.4799e-5
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_1=0.26523
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1=-0.12283
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_1=0.038525
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_2=0.050929
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_2=-0.033987
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_2=-6.2441e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_2=0.28227
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2=-0.12318
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_3=0.014657
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_3=-0.046178
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_3=4.5604e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_3=0.36575
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3=-0.14612
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4=-0.28
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_4=-4.0556e-7
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_4=-0.074414
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_4=0.00020273
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4=70000.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_4=1.6378e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5=-0.21656
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_5=-7.5152e-7
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_5=-0.05781
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_5=0.00030761
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5=-15180.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_5=4.8575e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_6=0.42387
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6=-0.16448
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_6=-0.053475
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_6=-0.040801
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_6=6.6904e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_7=-9.0e-12
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_7=0.42311
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7=-0.15062
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_7=0.0059558
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_7=-0.060009
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_7=0.00024431
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_8=0.35054
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8=-0.1508
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_8=0.0064044
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_8=-0.041595
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_8=8.2375e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_9=0.31431
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9=-0.15573
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_9=0.045814
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_9=-0.036237
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_9=6.5466e-5
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_10=0.00012837
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10=-0.13733
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_10=-0.035399
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_10=0.22183
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_10=0.084204
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_11=0.00023272
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11=57990.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11=-0.18157
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_11=-0.035319
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_12=-0.031044
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_12=0.059152
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_12=3.8701e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12=2640.7
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12=-0.15112
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_12=-2.0003e-6
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_13=-0.041096
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_13=0.31816
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_13=0.4
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_13=0.00017756
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13=-0.15
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_14=-0.039891
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_14=0.27573
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_14=0.051273
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_14=0.0002752
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14=-0.14408
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_15=-0.04584
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_15=0.32095
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_15=0.068491
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_15=0.00036886
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15=-0.18941
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_16=-0.046191
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_16=0.19162
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_16=0.10537
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_16=0.00022391
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16=-0.15862
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_17=-0.036588
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_17=0.18931
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_17=0.10003
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_17=0.0001803
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17=-0.14469
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_18=-0.036252
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_18=0.00019472
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18=80000.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18=-0.19865
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_19=-2.8735e-6
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_19=-0.036129
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_19=0.00079325
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_19=0.00034388
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19=1789.2
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19=-0.18947
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_20=-0.045969
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_20=0.36432
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_20=-0.08995
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_20=0.00027876
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20=-0.16549
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_21=0.00030084
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21=-0.16429
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_21=-9.0e-12
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_21=-0.059542
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_21=0.52752
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_21=-0.020825
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_22=0.38179
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_22=5.5575e-5
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_22=0.0002937
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22=-0.1684
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_22=-9.0e-12
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_22=-0.06861
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_23=-0.039682
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_23=0.16164
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_23=0.11227
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_23=0.00028783
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23=-0.1563
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_24=-0.039203
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_24=0.17776
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_24=0.10373
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_24=0.00030829
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24=-0.16924
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_25=-0.037386
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_25=0.00035668
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25=36375.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25=-0.1966
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_26=-0.040361
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_26=0.013843
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_26=0.00025252
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26=51375.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26=-0.15811
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_26=-1.9064e-6
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_27=-5.3555e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_27=4.9984e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_27=-0.075051
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_27=0.00077682
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27=-0.24948
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_28=-1.9408e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_28=2.0015e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_28=-0.031318
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_28=7.1455e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28=-0.07574
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_29=-2.4408e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_29=1.9709e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_29=-0.046346
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_29=0.0001927
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29=-0.13729
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_30=-2.2545e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_30=1.8478e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_30=-0.046449
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_30=0.00035799
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30=-0.14819
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_31=-1.9767e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_31=2.0771e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_31=-0.045925
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_31=0.00023018
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31=-0.12922
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_32=0.00013143
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32=77384.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32=-0.096134
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_32=-0.040413
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_33=0.00038874
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33=-16033.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33=-0.22536
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_33=-4.5931e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_33=2.1333e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_33=-0.063156
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_34=-0.059
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_34=0.00023588
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34=-0.14986
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_34=-4.2649e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_34=5.0e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_35=-0.028789
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_35=0.00018548
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35=-0.15
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_35=-3.1595e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_35=1.8164e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_36=-0.034578
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_36=0.00016852
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36=-0.15968
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_36=-4.7776e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_36=1.7566e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_37=1.9572e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_37=-0.024819
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_37=0.00021715
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37=-0.12769
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_37=-2.741e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_38=-0.054999
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_38=0.00027664
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38=80000.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38=-0.24782
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_39=-2.996e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_39=9.5527e-8
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_39=-0.070992
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_39=0.00080824
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39=15100.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39=-0.3
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_39=0.0
.include "sky130_fd_pr__pfet_01v8_lvt.pm3.spice"