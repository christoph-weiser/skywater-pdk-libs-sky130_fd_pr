* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8_lvt__toxe_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__overlap_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__ajunction_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__pjunction_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__lint_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__wint_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__dlc_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__dwc_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_37=0.0
.include "sky130_fd_pr__nfet_01v8_lvt.pm3.spice"