* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__special_nfet_pass_lvt__toxe_mult=1.052
.param sky130_fd_pr__special_nfet_pass_lvt__overlap_mult=0.98026
.param sky130_fd_pr__special_nfet_pass_lvt__ajunction_mult=1.1755
.param sky130_fd_pr__special_nfet_pass_lvt__pjunction_mult=1.0477
.param sky130_fd_pr__special_nfet_pass_lvt__rshn_mult=1.2
.param sky130_fd_pr__special_nfet_pass_lvt__lint_diff=-1.7325e-8
.param sky130_fd_pr__special_nfet_pass_lvt__wint_diff=3.2175e-8
.param sky130_fd_pr__special_nfet_pass_lvt__dlc_diff=-1.5633e-8
.param sky130_fd_pr__special_nfet_pass_lvt__dwc_diff=3.2175e-8
.param sky130_fd_pr__special_nfet_pass_lvt__u0_diff_0=5.0533e-3
.param sky130_fd_pr__special_nfet_pass_lvt__vsat_diff_0=5.6551e+4
.param sky130_fd_pr__special_nfet_pass_lvt__vth0_diff_0=1.6480e-1
.param sky130_fd_pr__special_nfet_pass_lvt__nfactor_diff_0=3.9755e-1
.param sky130_fd_pr__special_nfet_pass_lvt__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__ua_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__ub_diff_0=0.0
.include "sky130_fd_pr__special_nfet_pass_lvt.pm3.spice"