* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4_top c0 c1 m4 sub
xsky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4_0[0|0] c0 c1 m4 sub sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4
xsky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4_0[1|0] c0 c1 m4 sub sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4
xsky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4_0[0|1] c0 c1 m4 sub sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4
xsky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4_0[1|1] c0 c1 m4 sub sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4
.ends