* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__esd_nfet_01v8__toxe_mult=0.948
.param sky130_fd_pr__esd_nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__esd_nfet_01v8__overlap_mult=0.93416
.param sky130_fd_pr__esd_nfet_01v8__ajunction_mult=7.7394e-1
.param sky130_fd_pr__esd_nfet_01v8__pjunction_mult=7.9336e-1
.param sky130_fd_pr__esd_nfet_01v8__lint_diff=1.7325e-8
.param sky130_fd_pr__esd_nfet_01v8__wint_diff=-3.2175e-8
.param sky130_fd_pr__esd_nfet_01v8__dlc_diff=11.573e-9
.param sky130_fd_pr__esd_nfet_01v8__dwc_diff=-3.2175e-8
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_0=9.6384e-11
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_0=0.047703
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_0=-7.9399e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_0=-0.096312
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_0=-0.009208
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_0=-31425.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_0=-0.11707
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_1=5.9146e-11
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_1=0.023811
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_1=-5.5272e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_1=-0.095485
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_1=-0.0089632
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_1=-18149.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_1=-0.5032
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__esd_nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ags_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__ua_diff_2=5.8873e-11
.param sky130_fd_pr__esd_nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__a0_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__k2_diff_2=0.02267
.param sky130_fd_pr__esd_nfet_01v8__ub_diff_2=-8.0386e-19
.param sky130_fd_pr__esd_nfet_01v8__vth0_diff_2=-0.097368
.param sky130_fd_pr__esd_nfet_01v8__u0_diff_2=-0.0093619
.param sky130_fd_pr__esd_nfet_01v8__vsat_diff_2=-20000.0
.param sky130_fd_pr__esd_nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__nfactor_diff_2=-0.62007
.param sky130_fd_pr__esd_nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__esd_nfet_01v8__rdsw_diff_2=0.0
.include "sky130_fd_pr__esd_nfet_01v8.pm3.spice"