* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__special_nfet_pass_flash__tox_mult=1.0
.param sky130_fd_pr__special_nfet_pass_flash__ajunction_mult=9.9543e-1
.param sky130_fd_pr__special_nfet_pass_flash__pjunction_mult=1.0204e+0
.param sky130_fd_pr__special_nfet_pass_flash__overlap_mult=0.89805
.param sky130_fd_pr__special_nfet_pass_flash__lint_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__wint_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dwg_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__k3_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dvt0_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dvt0w_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__nlx_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cit_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cdsc_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cdscb_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__cdscd_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__kt2_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__kt1l_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dlc_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__dwc_diff=0.0
.param sky130_fd_pr__special_nfet_pass_flash__kt1_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_flash__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_flash__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_flash__u0_diff_0=0.0027584
.param sky130_fd_pr__special_nfet_pass_flash__vsat_diff_0=3855.4
.param sky130_fd_pr__special_nfet_pass_flash__vth0_diff_0=-0.15663
.param sky130_fd_pr__special_nfet_pass_flash__kt1_diff_1=3.8227e-2
.param sky130_fd_pr__special_nfet_pass_flash__nfactor_diff_1=1.4138e-1
.param sky130_fd_pr__special_nfet_pass_flash__voff_diff_1=0.0
.param sky130_fd_pr__special_nfet_pass_flash__k2_diff_1=0.0
.param sky130_fd_pr__special_nfet_pass_flash__u0_diff_1=1.2956e-3
.param sky130_fd_pr__special_nfet_pass_flash__vsat_diff_1=1.3679e+4
.param sky130_fd_pr__special_nfet_pass_flash__vth0_diff_1=-5.7093e-3
.param sky130_fd_pr__special_nfet_pass__tox_mult=1.0
.param sky130_fd_pr__special_nfet_pass__ajunction_mult=9.9543e-1
.param sky130_fd_pr__special_nfet_pass__pjunction_mult=1.0204e+0
.param sky130_fd_pr__special_nfet_pass__overlap_mult=0.9842
.param sky130_fd_pr__special_nfet_pass__lint_diff=0.0
.param sky130_fd_pr__special_nfet_pass__wint_diff=0.0
.param sky130_fd_pr__special_nfet_pass__k3_diff=0.0
.param sky130_fd_pr__special_nfet_pass__dvt0_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cit_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cdsc_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cdscb_diff=0.0
.param sky130_fd_pr__special_nfet_pass__cdscd_diff=0.0
.param sky130_fd_pr__special_nfet_pass__kt2_diff=0.0
.param sky130_fd_pr__special_nfet_pass__kt1l_diff=0.0
.param sky130_fd_pr__special_nfet_pass__dlc_diff=0.0
.param sky130_fd_pr__special_nfet_pass__dwc_diff=0.0
.param sky130_fd_pr__special_nfet_pass__kt1_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__nfactor_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__vsat_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__u0_diff_0=-0.0029226
.param sky130_fd_pr__special_nfet_pass__vth0_diff_0=0.027522
.param sky130_fd_pr__special_nfet_pass__rdsw_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__tox_mult=1.0
.param sky130_fd_pr__special_nfet_latch__ajunction_mult=9.9543e-1
.param sky130_fd_pr__special_nfet_latch__pjunction_mult=1.0204e+0
.param sky130_fd_pr__special_nfet_latch__overlap_mult=0.9842
.param sky130_fd_pr__special_nfet_latch__lint_diff=0.0
.param sky130_fd_pr__special_nfet_latch__wint_diff=0.0
.param sky130_fd_pr__special_nfet_latch__k3_diff=0.0
.param sky130_fd_pr__special_nfet_latch__dvt0_diff=0.0
.param sky130_fd_pr__special_nfet_latch__dvt1_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cit_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cdsc_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cdscb_diff=0.0
.param sky130_fd_pr__special_nfet_latch__cdscd_diff=0.0
.param sky130_fd_pr__special_nfet_latch__kt2_diff=0.0
.param sky130_fd_pr__special_nfet_latch__dlc_diff=0.0
.param sky130_fd_pr__special_nfet_latch__dwc_diff=0.0
.param sky130_fd_pr__special_nfet_latch__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__kt1_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__rdsw_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__u0_diff_0=0.00030368
.param sky130_fd_pr__special_nfet_latch__vth0_diff_0=0.020952
.param sky130_fd_pr__special_nfet_latch__vsat_diff_0=0.0
.param sky130_fd_pr__special_nfet_latch__nfactor_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__tox_mult=1.0
.param sky130_fd_pr__special_pfet_pass__ajunction_mult=9.9626e-1
.param sky130_fd_pr__special_pfet_pass__pjunction_mult=1.0009e+0
.param sky130_fd_pr__special_pfet_pass__overlap_mult=9.5435e-1
.param sky130_fd_pr__special_pfet_pass__lint_diff=0.0
.param sky130_fd_pr__special_pfet_pass__wint_diff=0.0
.param sky130_fd_pr__special_pfet_pass__k3_diff=0.0
.param sky130_fd_pr__special_pfet_pass__dvt0_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cit_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cdsc_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cdscb_diff=0.0
.param sky130_fd_pr__special_pfet_pass__cdscd_diff=0.0
.param sky130_fd_pr__special_pfet_pass__kt2_diff=0.0
.param sky130_fd_pr__special_pfet_pass__kt1l_diff=0.0
.param sky130_fd_pr__special_pfet_pass__dlc_diff=0.0
.param sky130_fd_pr__special_pfet_pass__dwc_diff=0.0
.param sky130_fd_pr__special_pfet_pass__voff_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__kt1_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__vsat_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__vth0_diff_0=0.0081943
.param sky130_fd_pr__special_pfet_pass__nfactor_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__k2_diff_0=0.0
.param sky130_fd_pr__special_pfet_pass__u0_diff_0=-0.00044468
.param sky130_fd_pr__special_pfet_pass__rdsw_diff_0=0.0
.include "../../../cells/special_nfet_latch/sky130_fd_pr__special_nfet_latch__mismatch.corner.spice"
.include "../../../cells/special_nfet_pass/sky130_fd_pr__special_nfet_pass__mismatch.corner.spice"
.include "../../../cells/special_nfet_pass_flash/sky130_fd_pr__special_nfet_pass_flash__mismatch.corner.spice"
.include "../../../cells/special_pfet_pass/sky130_fd_pr__special_pfet_pass__mismatch.corner.spice"
.include "../../../cells/special_nfet_pass_lvt/sky130_fd_pr__special_nfet_pass_lvt__tt.corner.spice"