* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff=0.0258
.param sky130_fd_pr__nfet_01v8_lvt__toxe_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__overlap_mult=9.2429e-1
.param sky130_fd_pr__nfet_01v8_lvt__ajunction_mult=1.0004e+0
.param sky130_fd_pr__nfet_01v8_lvt__pjunction_mult=8.9176e-1
.param sky130_fd_pr__nfet_01v8_lvt__lint_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__wint_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__dlc_diff=-1.3619e-9
.param sky130_fd_pr__nfet_01v8_lvt__dwc_diff=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_0=-0.070388
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_0=0.0081568
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_0=7.3798e-5
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_0=-0.12423
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_0=6.4377e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_0=2.3269e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0=0.89166
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0='-0.0042789+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_1=-0.064945
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_1=0.0073323
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_1=-0.14189
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_1=-0.00097736
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_1=3.5508e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_1=1.8212e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1=0.43195
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1='-0.0050888+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2='-0.0050675+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_2=0.0071155
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_2=0.0097539
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_2=0.022006
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_2=-0.0012946
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_2=-6.2443e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_2=1.6879e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2=0.87167
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3=1.5813
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3='-0.00024346+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_3=0.0025471
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_3=0.00016259
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_3=-1.4438e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3=-4935.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_3=1.6748e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4=1.6148
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4='-0.033357+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_4=0.0019871
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_4=-0.0014678
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_4=2.7231e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4=-6623.1
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_4=4.4948e-22
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_5=1.8383e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5=1.2444
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5='0.0058342+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_5=0.0054573
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_5=-0.0007973
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_5=-1.444e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5=-8609.7
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_6=1.2732e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6=1.2435
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6='-0.0052075+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_6=0.001201
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_6=-0.00049189
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_6=-5.5154e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6=2488.7
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_7=1.5266e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7=0.85875
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7='0.00035867+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_7=-0.05851
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_7=0.0048651
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_7=-0.074627
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_7=0.00064741
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_7=-1.2977e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_8=-0.080193
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_8=0.00048897
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_8=4.2479e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_8=1.7315e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8=0.40258
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8='-0.0059052+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_8=-0.0519
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_8=0.0029323
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_9=-0.011709
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_9=-0.00015331
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_9=-9.0975e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_9=1.0671e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9=0.51099
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9='-0.002435+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_9=0.0078569
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_9=0.0064203
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_10=3.9245e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_10=-3.2886e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_10=-0.0019115
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10=-778.01
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10='-0.039496+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10=1.3632
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_10=0.003079
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_11=0.0042111
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_11=1.1147e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_11=1.6097e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_11=0.00035625
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11=221.33
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11='-0.02476+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11=1.3783
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_12=0.0077253
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_12=1.6468e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_12=2.4517e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_12=-0.00021892
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12=1206.1
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12='-0.0039916+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12=1.0658
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_13=0.01115
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_13=-1.213e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_13=1.8252e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_13=0.00048299
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13=3587.4
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13='-0.0038667+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13=1.2498
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14=0.69102
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_14=0.0032333
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_14=-6.8844e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_14=1.7832e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_14=-0.062676
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_14=-0.090951
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_14=0.0009563
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14='-0.0067586+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15='-0.00026425+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15=0.63196
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_15=-0.0058846
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_15=-1.4976e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_15=1.8105e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_15=-0.0050262
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_15=-0.028351
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_15=0.00069251
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_16=-0.048053
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_16=0.00037829
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16='-0.0081622+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16=0.15108
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_16=0.009614
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_16=1.8675e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_16=1.4212e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_16=0.0077773
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_17=0.0004621
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17=3793.6
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17='-0.027423+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17=1.4437
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_17=0.002832
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_17=-1.0056e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_17=1.9308e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_18=-0.00039491
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18=-4510.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18='-0.011253+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18=1.3202
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_18=0.0049699
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_18=1.6514e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_18=1.2088e-19
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_19=1.6091e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_19=-0.0017408
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19=-5639.8
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19='-0.015458+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19=1.0129
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_19=0.0054353
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_19=3.4787e-12
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_20=-3.3561e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_20=2.4427e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_20=0.0015734
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20=5868.2
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20='-0.0087738+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20=1.04
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_20=0.0030478
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_21=-2.7372e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_21=2.0476e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_21=-0.0062986
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_21=-0.014108
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_21=0.0012828
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21='0.00055492+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21=0.75652
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_21=-0.0035982
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_22=0.0085737
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_22=-7.0145e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_22=1.5875e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_22=-0.024809
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_22=-0.065445
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_22=0.0006297
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22='-0.0047275+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22=0.4997
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_23=0.007571
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_23=-2.3602e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_23=2.0151e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_23=0.0034449
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_23=0.0091326
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_23=0.00087837
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23='-0.003912+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23=0.39236
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_24=0.0085689
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_24=6.3921e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_24=-1.368e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_24=-0.00323
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24=693.27
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24='-0.045182+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24=1.4575
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25=1.3049
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_25=0.006586
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_25=2.7798e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_25=1.0889e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_25=-0.00049693
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25=-1058.5
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25='-0.02251+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26='-0.012199+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26=1.0183
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_26=0.0067513
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_26=1.7984e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_26=2.6984e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_26=-0.00048946
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26=818.69
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_27=0.0011939
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27=-1097.6
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27='-0.0030064+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27=1.0842
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_27=0.0039291
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_27=-3.9545e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_27=2.1162e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_28=-0.0020626
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28='-0.0090378+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28=0.61174
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_28=8.0609e-8
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_28=2.2221e-9
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_28=0.00271
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_28=2.8232e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_28=2.5216e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_29=-0.00079351
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29=664.6
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29='-0.026469+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29=1.6428
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_29=0.0010093
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_29=7.1505e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_29=-3.5996e-20
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_30=4.6407e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_30=0.00050203
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30=-3707.1
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30='-0.044781+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30=1.5106
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_30=-0.00080889
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_30=4.4458e-12
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_31=1.5736e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_31=-2.585e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_31=-0.0019452
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31=-10041.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31='-0.02853+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31=1.9894
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_31=-0.0031204
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_32=1.2811e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_32=-1.4693e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_32=-0.0013308
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32=-1232.1
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32='-0.035332+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32=2.1559
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_32=-0.0040461
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_33=-0.0049622
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_33=8.2057e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_33=-1.3909e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_33=-0.0013932
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33=-1360.2
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33='-0.027481+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33=1.9686
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_34=0.004719
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_34=2.8047e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_34=-9.1484e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_34=-0.0023462
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34=252.46
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34='-0.026598+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34=1.4548
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_35=0.0022363
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_35=2.4112e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_35=-3.18e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_35=-0.0018653
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35=-3451.6
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35='-0.03725+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35=1.4139
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36=1.5691
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_36=0.0031583
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_36=-2.8757e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_36=2.2268e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_36=0.000508
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36=3914.9
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36='-0.025102+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37='-0.010883+sky130_fd_pr__nfet_01v8_lvt__vth0_correldiff'
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37=1.1341
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_37=0.0051762
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_37=2.2156e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_37=1.5682e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_37=-0.0017494
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37=-4160.7
.include "sky130_fd_pr__nfet_01v8_lvt.pm3.spice"