* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__rf_aura_blocking b_p d_n2 d_p d_p2 g g_n2 g_p g_p2 nwell s s_n2 s_p s_p2 vgnd vpwr
xsky130_fd_pr__rf_pfet_01v8_af02w3p00l0p15_0 d_p2 s_p2 g_p2 b_p subs sky130_fd_pr__rf_pfet_01v8_af02w3p00l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_0 d_n2 g_n2 s_n2 subs sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_0 d_p s_p g_p b_p subs sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_0 vpwr g s subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
.ends