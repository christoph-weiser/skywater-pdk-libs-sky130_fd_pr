* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre=0.0
.subckt sky130_fd_pr__nfet_01v8 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__nfet_01v8__model.0 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.5164001+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.026610291 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.68257 eta0=0.08 etab=-0.07 u0=0.0311586 ua=-7.5672677e-10 ub=1.58789e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.38376 ags=0.368846 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.1 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.5164001+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.026610291 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.68257 eta0=0.08 etab=-0.07 u0=0.0311586 ua=-7.5672677e-10 ub=1.58789e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.38376 ags=0.368846 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.2 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.169550527e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-4.439838262e-09 wvth0=-5.544600946e-08 pvth0=4.435897551e-13 k1=5.415455151e-01 lk1=-5.439186877e-09 wk1=-6.792616965e-08 pk1=5.434359163e-13 k2=-2.702810631e-02 lk2=3.342685843e-09 wk2=4.174444651e-08 pk2=-3.339718941e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.049995897e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.152187947e-09 wvoff=-2.687715773e-08 pvoff=2.150277708e-13 nfactor=2.684598982e+00 lnfactor=-1.623265138e-08 wnfactor=-2.027181371e-07 pnfactor=1.621824360e-12 eta0=0.08 etab=-0.07 u0=3.111987097e-02 lu0=3.098474224e-10 wu0=3.869465981e-09 pu0=-3.095724081e-14 ua=-7.563085878e-10 lua=-3.345620801e-18 wua=-4.178109914e-17 pua=3.342651295e-22 ub=1.582782613e-18 lub=4.086109167e-26 wub=5.102853621e-25 pub=-4.082482418e-30 uc=4.877028021e-11 luc=3.773942794e-18 wuc=4.713011049e-17 puc=-3.770593118e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.376602449e+00 la0=5.726320479e-08 wa0=7.151197875e-07 pa0=-5.721237912e-12 ags=3.702739278e-01 lags=-1.142398111e-08 wags=-1.426660449e-07 pags=1.141384142e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=1.950721142e-24 lb1=1.253031301e-30 wb1=1.564822438e-29 pb1=-1.251919135e-34 keta=-8.288268593e-03 lketa=-4.050849232e-09 wketa=-5.058819974e-08 pketa=4.047253779e-13 dwg=0.0 dwb=0.0 pclm=6.798847130e-02 lpclm=-3.333960644e-07 wpclm=-4.163548365e-06 ppclm=3.331001487e-11 pdiblc1=0.39 pdiblc2=3.074731630e-03 lpdiblc2=-1.018393736e-11 wpdiblc2=-1.271800128e-10 ppdiblc2=1.017489830e-15 pdiblcb=-0.025 drout=0.56 pscbe1=7.580428532e+08 lpscbe1=-2.695086297e+01 wpscbe1=-3.365703242e+02 ppscbe1=2.692694192e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.131868188e-01 lkt1=1.254611517e-09 wkt1=1.566795859e-08 pkt1=-1.253497949e-13 kt2=-4.539668283e-02 lkt2=6.667992640e-10 wkt2=8.327185837e-09 pkt2=-6.662074263e-14 at=140000.0 ute=-1.816358003e+00 lute=2.366518406e-08 wute=2.955377970e-07 pute=-2.364417931e-12 ua1=3.613815991e-10 lua1=1.171129310e-16 wua1=1.462540817e-15 pua1=-1.170089839e-20 ub1=-6.204561511e-19 lub1=-1.533182842e-25 wub1=-1.914683944e-24 pub1=1.531822019e-29 uc1=1.690943672e-11 luc1=-8.638211971e-18 wuc1=-1.078765384e-16 puc1=8.630544866e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.3 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.082895647e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.022550162e-08 wvth0=6.416054992e-08 pvth0=-3.488324862e-14 k1=5.303470136e-01 lk1=3.935919803e-08 wk1=1.368032768e-07 pk1=-2.755619188e-13 k2=-2.027781121e-02 lk2=-2.366113392e-08 wk2=-7.090368593e-08 pk2=1.166646810e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.377013124e-01 ldsub=8.920346908e-08 wdsub=2.227889570e-06 pdsub=-8.912429387e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.094468316e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.563851864e-08 wvoff=5.574887074e-08 pvoff=-1.155086498e-13 nfactor=2.656480338e+00 lnfactor=9.625292024e-08 wnfactor=-1.214596091e-07 pnfactor=1.296758476e-12 eta0=7.409084779e-02 leta0=2.363891931e-08 weta0=5.903907362e-07 peta0=-2.361793787e-12 etab=-6.483418875e-02 letab=-2.066526485e-08 wetab=-5.161226184e-07 petab=2.064692278e-12 u0=3.163793223e-02 lu0=-1.762600218e-09 wu0=4.183247760e-09 pu0=-3.221249061e-14 ua=-7.759969872e-10 lua=7.541567464e-17 wua=1.363035837e-15 pua=-5.285551897e-21 ub=1.676569356e-18 lub=-3.343225490e-25 wub=-1.992821733e-24 pub=5.930924676e-30 uc=5.886902198e-11 luc=-3.662497289e-17 wuc=-3.275870957e-16 puc=1.121956027e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.496166100e+00 la0=-4.210381484e-07 wa0=-1.606799823e-06 pa0=3.567348402e-12 ags=3.566728824e-01 lags=4.298551859e-08 wags=-7.037186914e-07 pags=3.385814099e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=4.528339301e-24 lb1=-9.058449182e-30 wb1=-3.129644877e-29 pb1=6.260513444e-35 keta=-1.648344570e-02 lketa=2.873306350e-08 wketa=8.740373469e-08 pketa=-1.472963146e-13 dwg=0.0 dwb=0.0 pclm=-6.199141083e-01 lpclm=2.418483224e-06 wpclm=8.534067672e-06 ppclm=-1.748541405e-11 pdiblc1=0.39 pdiblc2=3.181769776e-03 lpdiblc2=-4.383783715e-10 wpdiblc2=-1.253303843e-08 ppdiblc2=5.064577420e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.026020723e+08 lpscbe1=1.948339379e+02 wpscbe1=6.731406483e+02 ppscbe1=-1.346544495e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.112630179e-01 lkt1=-6.441344035e-09 wkt1=3.431256217e-08 pkt1=-1.999354992e-13 kt2=-4.402603391e-02 lkt2=-4.816332340e-09 wkt2=-1.655168082e-08 pkt2=3.290445163e-14 at=1.381373163e+05 lat=7.451463117e-03 wat=1.861030421e-01 pat=-7.444849348e-7 ute=-1.757396517e+00 lute=-2.122038146e-07 wute=-1.618132686e-06 pute=5.291012246e-12 ua1=6.250607809e-10 lua1=-9.377068951e-16 wua1=-5.199608359e-15 pua1=1.495030322e-20 ub1=-9.494904445e-19 lub1=1.162947542e-24 wub1=5.192390727e-24 pub1=-1.311285736e-29 uc1=-4.084632707e-13 luc1=6.064015931e-17 wuc1=1.706114446e-16 puc1=-2.510063339e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.4 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.252641416e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.730289106e-09 wvth0=-1.395901499e-07 pvth0=3.726978176e-13 k1=5.525319085e-01 lk1=-5.019266071e-09 wk1=-2.516422950e-07 pk1=5.014811071e-13 k2=-3.310977702e-02 lk2=2.007814991e-09 wk2=8.769929244e-08 pk2=-2.006032895e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.822943290e-01 wdsub=-2.227454103e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.030206999e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.783742727e-09 wvoff=1.370422496e-07 pvoff=-2.781271933e-13 nfactor=2.696066082e+00 lnfactor=1.706595406e-08 wnfactor=1.379166589e-06 pnfactor=-1.705080666e-12 eta0=8.605900740e-02 leta0=-3.020794611e-10 weta0=-6.053629548e-07 peta0=3.018113414e-14 etab=-7.515081076e-02 letab=-2.798703115e-11 wetab=5.146238999e-07 petab=2.796219042e-15 u0=3.048700444e-02 lu0=5.397053895e-10 wu0=1.503619859e-08 pu0=-5.392263578e-14 ua=-7.768031703e-10 lua=7.702835605e-17 wua=2.568023674e-15 pua=-7.695998722e-21 ub=1.548052532e-18 lub=-7.723865094e-26 wub=-2.885689612e-24 pub=7.717009546e-30 uc=3.956086411e-11 luc=1.998892326e-18 wuc=3.331176577e-16 puc=-1.997118149e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.150917279e+04 lvsat=-3.018935661e-03 wvsat=-1.507833276e-01 pvsat=3.016256114e-7 a0=1.273571673e+00 la0=2.423774059e-08 wa0=1.387100453e-06 pa0=-2.421622766e-12 ags=4.017765750e-01 lags=-4.723950215e-08 wags=-1.370559940e-06 pags=4.719757332e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.947922130e-03 lketa=9.658287975e-09 wketa=4.961614388e-07 pketa=-9.649715472e-13 dwg=0.0 dwb=0.0 pclm=5.766408394e-01 lpclm=2.490547562e-08 wpclm=1.036994827e-06 ppclm=-2.488337002e-12 pdiblc1=4.135789662e-01 lpdiblc1=-4.716715180e-08 wpdiblc1=-2.355803799e-06 ppdiblc1=4.712528718e-12 pdiblc2=2.903068620e-03 lpdiblc2=1.191329119e-10 wpdiblc2=1.873509434e-08 ppdiblc2=-1.190271719e-14 pdiblcb=-2.315565645e-02 lpdiblcb=-3.689408231e-09 wpdiblcb=-1.842706544e-07 ppdiblcb=3.686133586e-13 drout=5.376969539e-01 ldrout=4.461481272e-08 wdrout=2.228325038e-06 pdrout=-4.457521351e-12 pscbe1=7.599344035e+08 lpscbe1=8.014685859e+01 wpscbe1=4.003003505e+03 ppscbe1=-8.007572184e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.240365012e-07 lalpha0=-3.881488707e-13 walpha0=-1.938642783e-11 palpha0=3.878043575e-17 alpha1=8.525276786e-01 lalpha1=-5.056345442e-09 walpha1=-2.525435043e-07 palpha1=5.051857531e-13 beta0=1.406608015e+01 lbeta0=-4.122408695e-07 wbeta0=-2.058972335e-05 pbeta0=4.118749728e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.106699830e-01 lkt1=-7.627645815e-09 wkt1=-4.466049515e-07 pkt1=7.620875669e-13 kt2=-4.494226573e-02 lkt2=-2.983510458e-09 wkt2=-1.491166563e-07 pkt2=2.980862354e-13 at=1.380281286e+05 lat=7.669881171e-03 wat=1.970121189e-01 pat=-7.663073538e-7 ute=-1.801915273e+00 lute=-1.231488964e-07 wute=-5.123920776e-06 pute=1.230395919e-11 ua1=2.840854611e-10 lua1=-2.556229341e-16 wua1=-1.049322426e-14 pua1=2.553960483e-20 ub1=-4.352212600e-19 lub1=1.342080935e-25 wub1=5.340381770e-24 pub1=-1.340889731e-29 uc1=3.135027395e-11 luc1=-2.889732799e-18 wuc1=-9.919737126e-17 puc1=2.887167930e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.5 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.167505171e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.786664210e-09 wvth0=8.181352179e-08 pvth0=1.512075771e-13 k1=5.403718237e-01 lk1=7.145573309e-09 wk1=9.760905180e-07 pk1=-7.267317495e-13 k2=-2.642553407e-02 lk2=-4.679041500e-09 wk2=-4.106816328e-07 pk2=2.979725027e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=9.149182842e-01 ldsub=-3.327540112e-07 wdsub=-5.463514810e-06 pdsub=3.237326006e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.009638102e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.260487701e-10 wvoff=-4.160901059e-08 pvoff=-9.940608042e-14 nfactor=2.651631826e+00 lnfactor=6.151758342e-08 wnfactor=-1.275597735e-06 pnfactor=9.507216707e-13 eta0=2.074861233e-01 leta0=-1.217766734e-07 weta0=-4.788141797e-06 peta0=4.214595442e-12 etab=-1.499012846e-01 letab=7.475171430e-08 wetab=1.033844291e-06 petab=-5.166271874e-13 u0=3.263025303e-02 lu0=-1.604381218e-09 wu0=-3.857549189e-08 pu0=-2.899831220e-16 ua=-5.269283583e-10 lua=-1.729441569e-16 wua=-5.170155120e-15 pua=4.520570007e-23 ub=1.334918308e-18 lub=1.359789082e-25 wub=5.318206731e-24 pub=-4.900945202e-31 uc=9.405668330e-12 luc=3.216587879e-17 wuc=2.043946234e-16 puc=-7.093844997e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.973799759e+04 lvsat=-1.247067935e-03 wvsat=2.617698615e-02 pvsat=1.245961062e-7 a0=1.298398683e+00 la0=-5.989771743e-10 wa0=-3.470644325e-06 pa0=2.438021390e-12 ags=2.419393853e-01 lags=1.126601839e-07 wags=1.282167580e-06 pags=2.065992595e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.555209912e-03 lketa=-8.489507921e-10 wketa=-7.386578190e-07 pketa=2.703305250e-13 dwg=0.0 dwb=0.0 pclm=6.422792070e-01 lpclm=-4.075855658e-08 wpclm=-2.734312189e-06 ppclm=1.284444595e-12 pdiblc1=3.882093194e-01 lpdiblc1=-2.178758547e-08 wpdiblc1=1.789091215e-07 ppdiblc1=2.176824724e-12 pdiblc2=1.127247562e-03 lpdiblc2=1.895648316e-09 wpdiblc2=2.398714120e-08 ppdiblc2=-1.715681759e-14 pdiblcb=-2.868868709e-02 lpdiblcb=1.845785823e-09 wpdiblcb=3.685413088e-07 ppdiblcb=-1.844147540e-13 drout=6.000509517e-01 ldrout=-1.776356547e-08 wdrout=-4.001540324e-06 pdrout=1.774779888e-12 pscbe1=8.623427798e+08 lpscbe1=-2.230155932e+01 wpscbe1=-6.228744556e+03 ppscbe1=2.228176491e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=8.593108523e-08 lalpha0=-2.499894555e-13 walpha0=-5.588144192e-12 palpha0=2.497675698e-17 alpha1=8.449446429e-01 lalpha1=2.529655204e-09 walpha1=5.050870086e-07 palpha1=-2.527409933e-13 beta0=1.381524008e+01 lbeta0=-1.613027201e-07 wbeta0=4.472019687e-06 pbeta0=1.611595510e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.090922339e-01 lkt1=-9.206011784e-09 wkt1=2.796662331e-07 pkt1=3.553241023e-14 kt2=-4.863049774e-02 lkt2=7.061636498e-10 wkt2=2.207618376e-07 pkt2=-7.193688096e-14 at=1.718992706e+05 lat=-2.621450440e-02 wat=-6.813620641e-01 pat=1.124102735e-7 ute=-2.113891966e+00 lute=1.889497800e-07 wute=1.221752792e-05 pute=-5.044270011e-12 ua1=-3.811741320e-10 lua1=4.098967755e-16 wua1=2.534894290e-14 pua1=-1.031657662e-20 ub1=-8.376487019e-20 lub1=-2.173857157e-25 wub1=-1.142201320e-23 pub1=3.360051755e-30 uc1=1.675069851e-11 luc1=1.171555108e-17 wuc1=7.516671442e-16 puc1=-5.624804104e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.6 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.227182158e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.800481472e-09 wvth0=7.434879268e-07 pvth0=-1.798883401e-13 k1=5.751953467e-01 lk1=-1.027980420e-08 wk1=-2.528768193e-06 pk1=1.027068006e-12 k2=-4.206457837e-02 lk2=3.146595520e-09 wk2=8.130669341e-07 pk2=-3.143802665e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.620200156e-01 ldsub=-6.049593613e-09 wdsub=-2.018222635e-07 pdsub=6.044224115e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.001123163e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.999688846e-10 wvoff=-1.803721310e-07 pvoff=-2.997026382e-14 nfactor=2.794368815e+00 lnfactor=-9.906720777e-09 wnfactor=-1.353678888e-06 pnfactor=9.897927770e-13 eta0=-3.587691354e-02 weta0=3.634462612e-6 etab=-5.576476861e-04 letab=2.150245380e-11 wetab=5.690606260e-09 petab=-2.148336865e-15 u0=2.884172015e-02 lu0=2.913665383e-10 wu0=1.902108677e-08 pu0=-2.911079271e-14 ua=-9.107021033e-10 lua=1.909277112e-17 wua=-1.267630543e-15 pua=-1.907582476e-21 ub=1.625779571e-18 lub=-9.565450053e-27 wub=2.428885150e-24 pub=9.556959951e-31 uc=7.382403576e-11 luc=-6.849250921e-20 wuc=4.895293557e-17 puc=6.843171663e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.033205551e+04 lvsat=-1.544329172e-03 wvsat=-3.317607853e-02 pvsat=1.542958456e-7 a0=1.297201665e+00 wa0=1.401588370e-6 ags=3.754990731e-01 lags=4.582811817e-08 wags=1.456125693e-05 pags=-4.578744205e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=9.873100969e-04 lketa=4.360031644e-10 wketa=-1.113640774e-07 pketa=-4.356161767e-14 dwg=0.0 dwb=0.0 pclm=5.515509861e-01 lpclm=4.641028587e-09 wpclm=7.592269146e-07 ppclm=-4.636909303e-13 pdiblc1=2.790320437e-01 lpdiblc1=3.284374068e-08 wpdiblc1=1.108694633e-05 ppdiblc1=-3.281458923e-12 pdiblc2=4.849674909e-03 lpdiblc2=3.297917298e-11 wpdiblc2=-3.714850765e-09 ppdiblc2=-3.294990132e-15 pdiblcb=-3.988613158e-02 lpdiblcb=7.448886265e-09 wpdiblcb=1.487291894e-06 ppdiblcb=-7.442274783e-13 drout=6.018597706e-01 ldrout=-1.866868219e-08 wdrout=-4.182261671e-06 pdrout=1.865211224e-12 pscbe1=8.355768263e+08 lpscbe1=-8.908117125e+00 wpscbe1=-3.554524907e+03 ppscbe1=8.900210459e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.637441582e-07 lalpha0=1.251412893e-13 walpha0=6.931284048e-11 palpha0=-1.250302163e-17 alpha1=0.85 beta0=1.351722554e+01 lbeta0=-1.217892904e-08 wbeta0=3.424702199e-05 pbeta0=1.216811927e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.285997835e-01 lkt1=5.553904497e-10 wkt1=4.615683054e-07 pkt1=-5.548974962e-14 kt2=-4.750756286e-02 lkt2=1.442571426e-10 wkt2=1.058037935e-07 pkt2=-1.441291029e-14 at=1.174641194e+05 lat=1.024355308e-03 wat=-2.521879090e-01 pat=-1.023446111e-7 ute=-1.694739682e+00 lute=-2.079025088e-08 wute=-2.014242434e-06 pute=2.077179787e-12 ua1=4.631243163e-10 lua1=-1.258256929e-17 wua1=2.219596551e-15 pua1=1.257140126e-21 ub1=-4.860441619e-19 lub1=-1.608877868e-26 wub1=-7.919548334e-24 pub1=1.607449860e-30 uc1=4.788836180e-11 luc1=-3.865455391e-18 wuc1=-1.144215994e-15 puc1=3.862024490e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.7 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.217879014e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.033423839e-09 wvth0=8.364367992e-07 pvth0=-2.031619012e-13 k1=5.580741000e-01 lk1=-5.992798130e-09 wk1=-8.181631732e-07 pk1=5.987479042e-13 k2=-3.813298494e-02 lk2=2.162159909e-09 wk2=4.202565515e-07 pk2=-2.160240819e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.074114547e-01 ldsub=7.623898551e-09 wdsub=5.254186876e-06 pdsub=-7.617131731e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.013136585e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.007741479e-10 wvoff=-6.034454434e-08 pvoff=-6.002409128e-14 nfactor=2.779488868e+00 lnfactor=-6.180916116e-09 wnfactor=1.329950388e-07 pnfactor=6.175430059e-13 eta0=-1.237830042e-01 leta0=2.201089394e-08 weta0=1.241726931e-05 peta0=-2.199135751e-12 etab=-5.732090360e-03 letab=1.317136329e-09 wetab=5.226756005e-07 petab=-1.315967266e-13 u0=3.284169641e-02 lu0=-7.101915170e-10 wu0=-3.806215092e-07 pu0=7.095611652e-14 ua=-5.723411799e-10 lua=-6.562975886e-17 wua=-3.507369065e-14 pua=6.557150720e-21 ub=1.418298767e-18 lub=4.238587584e-26 wub=2.315854993e-23 pub=-4.234825498e-30 uc=7.389731697e-11 luc=-8.684146528e-20 wuc=4.163131861e-17 puc=8.676438653e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.493865736e+04 lvsat=-1.938708140e-04 wvsat=5.056850298e-01 pvsat=1.936987381e-8 a0=1.297201665e+00 wa0=1.401588370e-6 ags=7.941716087e-01 lags=-5.900371670e-08 wags=-2.726883609e-05 pags=5.895134618e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.597134530e-03 lketa=3.291761466e-11 wketa=-2.722036359e-07 pketa=-3.288839764e-15 dwg=0.0 dwb=0.0 pclm=5.460401978e-01 lpclm=6.020880387e-09 wpclm=1.309816620e-06 ppclm=-6.015536374e-13 pdiblc1=4.593656043e-01 lpdiblc1=-1.231015988e-08 wpdiblc1=-6.930403679e-06 ppdiblc1=1.229923363e-12 pdiblc2=6.185918179e-03 lpdiblc2=-3.016041156e-10 wpdiblc2=-1.372205755e-07 ppdiblc2=3.013364178e-14 pdiblcb=1.641448547e-02 lpdiblcb=-6.648281538e-09 wpdiblcb=-4.137772680e-06 ppdiblcb=6.642380656e-13 drout=4.730856358e-01 ldrout=1.357520219e-08 wdrout=8.683722070e-06 pdrout=-1.356315311e-12 pscbe1=7.992141395e+08 lpscbe1=1.967724026e-01 wpscbe1=7.851630106e+01 ppscbe1=-1.965977514e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.676681667e-07 lalpha0=1.261238257e-13 walpha0=6.970489304e-11 palpha0=-1.260118807e-17 alpha1=9.153238386e-01 lalpha1=-1.635650127e-08 walpha1=-6.526585848e-06 palpha1=1.634198357e-12 beta0=1.267822682e+01 lbeta0=1.978988002e-07 wbeta0=1.180724264e-04 pbeta0=-1.977231492e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.201512214e-01 lkt1=-1.560053457e-09 wkt1=-3.825380247e-07 pkt1=1.558668785e-13 kt2=-4.620558524e-02 lkt2=-1.817463356e-10 wkt2=-2.427840760e-08 pkt2=1.815850212e-14 at=1.234782819e+05 lat=-4.815368361e-04 wat=-8.530703467e-01 pat=4.811094336e-8 ute=-1.960769993e+00 lute=4.582134483e-08 wute=2.456517639e-05 pute=-4.578067472e-12 ua1=2.689415591e-11 lua1=9.664553680e-17 wua1=4.580389367e-14 pua1=-9.655975615e-21 ub1=-2.277319808e-19 lub1=-8.076782403e-26 wub1=-3.372783918e-23 pub1=8.069613612e-30 uc1=4.041130723e-11 luc1=-1.993268220e-18 wuc1=-3.971741856e-16 puc1=1.991499035e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.8 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.265882882e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.167477261e-09 wvth0=3.568241907e-07 pvth0=-1.166441032e-13 k1=5.308143895e-01 lk1=-1.075391689e-09 wk1=1.905388362e-06 pk1=1.074437193e-13 k2=-3.070339202e-02 lk2=8.219282118e-10 wk2=-3.220433053e-07 pk2=-8.211986848e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.226984096e-01 ldsub=4.866269467e-09 wdsub=3.726848225e-06 pdsub=-4.861950264e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=3.388280476e-03 lcdscd=3.628961577e-10 wcdscd=2.009934300e-07 pcdscd=-3.625740583e-14 cit=0.0 voff='-1.214533238e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.233788507e-09 wvoff=1.951834427e-06 pvoff=-4.230030681e-13 nfactor=1.992446753e+00 lnfactor=1.357943982e-07 wnfactor=7.876735031e-05 pnfactor=-1.356738698e-11 eta0=-1.301640020e-02 leta0=2.029595483e-09 weta0=1.350440331e-06 peta0=-2.027794055e-13 etab=-3.731961242e-03 letab=9.563310376e-10 wetab=3.228402161e-07 petab=-9.554822173e-14 u0=2.448748741e-02 lu0=7.968325985e-10 wu0=4.540578878e-07 pu0=-7.961253458e-14 ua=-1.520016895e-09 lua=1.053224110e-16 wua=5.960976703e-14 pua=-1.052289289e-20 ub=2.170143346e-18 lub=-9.324011946e-26 wub=-5.195917567e-23 pub=9.315736139e-30 uc=6.102110797e-11 luc=2.235910752e-18 wuc=1.328109352e-15 puc=-2.233926203e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.925236073e+04 lvsat=-9.720240787e-04 wvsat=7.469756841e-02 pvsat=9.711613296e-8 a0=1.297201665e+00 wa0=1.401588370e-6 ags=4.670836902e-01 wags=5.410924083e-6 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.578400295e-02 lketa=-4.149784766e-09 wketa=-2.588832458e-06 pketa=4.146101501e-13 dwg=0.0 dwb=0.0 pclm=5.358521201e-01 lpclm=7.858717904e-09 wpclm=2.327720113e-06 ppclm=-7.851742663e-13 pdiblc1=3.955332388e-01 lpdiblc1=-7.953756376e-10 wpdiblc1=-5.528327618e-07 ppdiblc1=7.946696781e-14 pdiblc2=4.783093782e-03 lpdiblc2=-4.854721977e-11 wpdiblc2=2.937352361e-09 ppdiblc2=4.850413023e-15 pdiblcb=1.172724263e-02 lpdiblcb=-5.802745115e-09 wpdiblcb=-3.669464427e-06 ppdiblcb=5.797594714e-13 drout=4.811642345e-01 ldrout=1.211789570e-08 wdrout=7.876579247e-06 pdrout=-1.210714010e-12 pscbe1=7.983077928e+08 lpscbe1=3.602691928e-01 wpscbe1=1.690705270e+02 ppscbe1=-3.599494250e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.902558023e-08 lalpha0=-1.357366036e-15 walpha0=-9.017569302e-13 palpha0=1.356161265e-19 alpha1=6.975777099e-01 lalpha1=2.292294063e-08 walpha1=1.522870031e-05 palpha1=-2.290259469e-12 beta0=1.335058513e+01 lbeta0=7.661141107e-08 wbeta0=5.089627193e-05 pbeta0=-7.654341232e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.125161885e-01 lkt1=-2.937344671e-09 wkt1=-1.145363641e-06 pkt1=2.934737543e-13 kt2=-4.470679961e-02 lkt2=-4.521137749e-10 wkt2=-1.740239417e-07 pkt2=4.517124877e-14 at=1.196028009e+05 lat=2.175650501e-04 wat=-4.658662305e-01 pat=-2.173719438e-8 ute=-1.027076231e+00 lute=-1.226086066e-07 wute=-6.872132702e-05 pute=1.224997816e-11 ua1=1.509264701e-09 lua1=-1.707607682e-16 wua1=-1.023015886e-13 pua1=1.706092044e-20 ub1=-1.217957253e-18 lub1=9.785990313e-26 wub1=6.520679767e-23 pub1=-9.777304464e-30 uc1=3.948670632e-11 luc1=-1.826478539e-18 wuc1=-3.047961609e-16 puc1=1.824857393e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.9 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.183061289e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.906036344e-07 wvth0=-1.317302693e-08 pvth0=1.317307844e-12 k1=5.418096583e-01 lk1=-9.440119709e-08 wk1=-6.524269672e-09 pk1=6.524295182e-13 k2=-2.732440569e-02 lk2=7.141174787e-08 wk2=4.935419414e-09 pk2=-4.935438712e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.045392417e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.293611037e-08 wvoff=-5.040771383e-09 pvoff=5.040791093e-13 nfactor=2.602103866e+00 lnfactor=8.046644882e-06 wnfactor=5.561209263e-07 pnfactor=-5.561231007e-11 eta0=0.08 etab=-0.07 u0=3.108707864e-02 lu0=7.152163949e-09 wu0=4.943014260e-10 pu0=-4.943033587e-14 ua=-7.350589596e-10 lua=-2.166789508e-15 wua=-1.497514810e-16 pua=1.497520665e-20 ub=1.548267781e-18 lub=3.962237436e-24 wub=2.738387471e-25 pub=-2.738398178e-29 uc=4.773237748e-11 luc=1.509628425e-16 wuc=1.043336658e-17 puc=-1.043340737e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.392893247e+00 la0=-9.133282667e-07 wa0=-6.312207996e-08 pa0=6.312232676e-12 ags=3.689872010e-01 lags=-1.412015200e-08 wags=-9.758740600e-10 pags=9.758778756e-14 a1=0.0 a2=0.42385546 b0=0.0 b1=8.136085451e-25 lb1=1.293738913e-28 wb1=8.941307755e-30 pb1=-8.941342715e-34 keta=-7.193719169e-03 lketa=-1.600887090e-07 wketa=-1.106407483e-08 pketa=1.106411809e-12 dwg=0.0 dwb=0.0 pclm=5.735933976e-02 lpclm=-3.104346114e-06 wpclm=-2.145480335e-07 ppclm=2.145488724e-11 pdiblc1=0.39 pdiblc2=3.147270094e-03 lpdiblc2=-7.381168258e-09 wpdiblc2=-5.101284061e-10 ppdiblc2=5.101304007e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.177508068e+08 lpscbe1=3.692349762e+03 wpscbe1=2.551862297e+02 ppscbe1=-2.551872275e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.200102392e-01 lkt1=6.980266446e-07 wkt1=4.824212201e-08 pkt1=-4.824231063e-12 kt2=-4.543376669e-02 lkt2=1.204301625e-08 wkt2=8.323187428e-10 pkt2=-8.323219972e-14 at=140000.0 ute=-1.856558383e+00 lute=4.315855155e-06 wute=2.982780279e-07 pute=-2.982791942e-11 ua1=3.042407949e-10 lua1=7.177948574e-15 wua1=4.960834569e-16 pua1=-4.960853966e-20 ub1=-5.525849512e-19 lub1=-8.703538910e-24 wub1=-6.015202847e-25 pub1=6.015226366e-29 uc1=1.656470333e-11 luc1=-7.349932026e-17 wuc1=-5.079696030e-18 puc1=5.079715891e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.10 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.087761335e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=5.269107761e-8 k1=5.370896907e-01 wk1=2.609656850e-8 k2=-2.375388810e-02 wk2=-1.974129171e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.081859760e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=2.016269135e-8 nfactor=3.004428244e+00 wnfactor=-2.224440217e-6 eta0=0.08 etab=-0.07 u0=3.144467985e-02 wu0=-1.977167050e-9 ua=-8.433963170e-10 wua=5.989942136e-16 ub=1.746375779e-18 wub=-1.095333575e-24 uc=5.528037204e-11 wuc=-4.173265045e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.347227726e+00 wa0=2.524833838e-7 ags=3.682812072e-01 wags=3.903419928e-9 a1=0.0 a2=0.42385546 b0=0.0 b1=7.282176652e-24 wb1=-3.576453182e-29 keta=-1.519799814e-02 wketa=4.425543414e-8 dwg=0.0 dwb=0.0 pclm=-9.785493149e-02 wpclm=8.581753569e-7 pdiblc1=0.39 pdiblc2=2.778218896e-03 wpdiblc2=2.040473733e-9 pdiblcb=-0.025 drout=0.56 pscbe1=9.023646856e+08 wpscbe1=-1.020724964e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.851095892e-01 wkt1=-1.929647156e-7 kt2=-4.483162765e-02 wkt2=-3.329209885e-9 at=140000.0 ute=-1.640769844e+00 wute=-1.193088787e-6 ua1=6.631312073e-10 wua1=-1.984295035e-15 ub1=-9.877533892e-19 wub1=2.406034101e-24 uc1=1.288980916e-11 wuc1=2.031838689e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.11 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.945801811e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.135731696e-07 wvth0=9.919214254e-08 pvth0=-3.720267014e-13 k1=5.247002949e-01 lk1=9.912001029e-08 wk1=4.849522359e-08 pk1=-1.791979986e-13 k2=-1.341469649e-02 lk2=-8.271757551e-08 wk2=-5.234112323e-08 pk2=2.608113986e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.176212750e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.548608176e-08 wvoff=6.035436443e-08 pvoff=-3.215490996e-13 nfactor=3.334011302e+00 lnfactor=-2.636793325e-06 wnfactor=-4.690963835e-06 pnfactor=1.973315335e-11 eta0=0.08 etab=-0.07 u0=3.236097882e-02 lu0=-7.330750100e-09 wu0=-4.708130787e-09 pu0=2.184877770e-14 ua=-8.816945241e-10 lua=3.064006308e-16 wua=8.247914495e-16 pua=-1.806466174e-21 ub=1.939418182e-18 lub=-1.544414704e-24 wub=-1.954509363e-24 pub=6.873742243e-30 uc=1.750887724e-10 luc=-9.585140477e-16 wuc=-8.258875579e-16 puc=6.273545864e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.744134619e+00 la0=-3.175410335e-06 wa0=-1.824983983e-06 pa0=1.662055123e-11 ags=4.446122939e-01 lags=-6.106785396e-07 wags=-6.564364828e-07 pags=5.282977415e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=1.456506514e-23 lb1=-5.826595548e-29 wb1=-7.153255963e-29 pb1=2.861582077e-34 keta=-2.846204951e-02 lketa=1.061175972e-07 wketa=8.883768220e-08 pketa=-3.566754161e-13 dwg=0.0 dwb=0.0 pclm=-1.020401365e+00 lpclm=7.380732182e-06 wpclm=3.358577183e-06 ppclm=-2.000419226e-11 pdiblc1=0.39 pdiblc2=2.817055066e-03 lpdiblc2=-3.107045406e-10 wpdiblc2=1.653685082e-09 ppdiblc2=3.094460445e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.002114750e+09 lpscbe1=-7.980395141e+02 wpscbe1=-2.023410265e+03 ppscbe1=8.021874464e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.599879651e-01 lkt1=-2.009828159e-07 wkt1=-3.520021936e-07 pkt1=1.272362008e-12 kt2=-3.218308448e-02 lkt2=-1.011932910e-07 wkt2=-8.299519008e-08 pkt2=6.373589910e-13 at=140000.0 ute=-1.122318637e+00 lute=-4.147812367e-06 wute=-4.501136221e-06 pute=2.646567292e-11 ua1=1.914829100e-09 lua1=-1.001407255e-14 wua1=-9.273710794e-15 pua1=5.831817624e-20 ub1=-2.188679232e-18 lub1=9.607876306e-24 wub1=8.923685280e-24 pub1=-5.214375783e-29 uc1=-2.772335591e-11 luc1=3.249212003e-16 wuc1=2.005914926e-16 puc1=-1.442255333e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.12 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.209634013e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.029972927e-09 wvth0=-2.343140173e-08 pvth0=1.185154215e-13 k1=5.756201135e-01 lk1=-1.045791735e-07 wk1=-1.760900728e-07 pk1=7.192310000e-13 k2=-4.238690165e-02 lk2=3.318257327e-08 wk2=8.189758849e-08 pk2=-2.761959356e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.871463510e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.015178051e-08 wvoff=-8.753635636e-08 pvoff=2.700716089e-13 nfactor=2.578836738e+00 lnfactor=3.842002027e-07 wnfactor=4.151540995e-07 pnfactor=-6.933148763e-13 eta0=1.595155422e-01 leta0=-3.180932596e-7 etab=-1.395111990e-01 letab=2.780719748e-07 wetab=-1.172884486e-11 petab=4.691996542e-17 u0=3.190674932e-02 lu0=-5.513654492e-09 wu0=2.325387804e-09 pu0=-6.288046772e-15 ua=-4.012728211e-10 lua=-1.615474026e-15 wua=-1.226773558e-15 pua=6.400596019e-21 ub=1.016314898e-18 lub=2.148359367e-24 wub=2.570356607e-24 pub=-1.122749086e-29 uc=-2.094599961e-10 luc=5.798313848e-16 wuc=1.526899684e-15 puc=-3.138523043e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=4.829221617e-01 la0=1.869932630e-06 wa0=5.395974240e-06 pa0=-1.226610506e-11 ags=1.007210087e-01 lags=7.650210627e-07 wags=1.065226648e-06 pags=-1.604348279e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.666402628e-05 lketa=-7.635062953e-09 wketa=-2.633306598e-08 pketa=1.040526084e-13 dwg=0.0 dwb=0.0 pclm=8.328770938e-01 lpclm=-3.310628388e-08 wpclm=-1.506523901e-06 ppclm=-5.418856722e-13 pdiblc1=0.39 pdiblc2=1.313149826e-03 lpdiblc2=5.705504444e-09 wpdiblc2=3.814462430e-10 ppdiblc2=8.183913246e-15 pdiblcb=-0.025 drout=0.56 pscbe1=8.052492556e+08 lpscbe1=-1.050056369e+01 wpscbe1=-3.627887587e+01 ppscbe1=7.257193679e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.046290832e-01 lkt1=-2.240088868e-08 wkt1=-1.153616624e-08 pkt1=-8.963522397e-14 kt2=-5.804798575e-02 lkt2=2.276427313e-09 wkt2=8.035742164e-08 pkt2=-1.611532678e-14 at=1.680859036e+05 lat=-1.123545958e-01 wat=-2.087889194e-02 pat=8.352373143e-8 ute=-2.533283117e+00 lute=1.496597241e-06 wute=3.744207372e-06 pute=-6.518925380e-12 ua1=-1.720721890e-09 lua1=4.529552908e-15 wua1=1.101266336e-14 pua1=-2.283525236e-20 ub1=1.239220991e-18 lub1=-4.105064897e-24 wub1=-9.934323674e-24 pub1=2.329565147e-29 uc1=6.704513814e-11 luc1=-5.418983040e-17 wuc1=-2.955767185e-16 puc1=5.426115138e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.13 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.009590040e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.804658922e-08 wvth0=2.838853748e-08 pvth0=1.485528149e-14 k1=4.326433527e-01 lk1=1.814302520e-07 wk1=5.769365271e-07 pk1=-7.871166332e-13 k2=1.002041037e-02 lk2=-7.165254202e-08 wk2=-2.103838701e-07 pk2=3.084812637e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.146671521e+00 ldsub=-1.773689731e-06 wdsub=-6.128001457e-06 pdsub=1.225839896e-11 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.037666527e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.004185994e-08 wvoff=1.421977098e-07 pvoff=-1.894863494e-13 nfactor=2.844007348e+00 lnfactor=-1.462446987e-07 wnfactor=3.567086993e-07 pnfactor=-5.764012239e-13 eta0=-6.536868951e-03 leta0=1.407648932e-08 weta0=3.458955489e-08 peta0=-6.919263430e-14 etab=-9.720590370e-04 letab=9.395261037e-10 wetab=1.956595516e-09 petab=-3.890498372e-15 u0=3.281190827e-02 lu0=-7.324326295e-09 wu0=-1.031774403e-09 pu0=4.275902925e-16 ua=-9.154920735e-10 lua=-5.868344616e-16 wua=3.526536247e-15 pua=-3.107882135e-21 ub=1.951553603e-18 lub=2.775162797e-25 wub=-5.674383160e-24 pub=5.265212370e-30 uc=7.458568807e-11 luc=1.162895455e-17 wuc=9.105262328e-17 puc=-2.662675054e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.932552128e+04 lvsat=1.213726812e-01 wvsat=2.789829365e-01 pvsat=-5.580749553e-7 a0=2.274545452e+00 la0=-1.714014475e-06 wa0=-5.530871569e-06 pa0=9.591858953e-12 ags=9.550908884e-01 lags=-9.440527552e-07 wags=-5.194649062e-06 pags=1.091785075e-11 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.292897922e-02 lketa=-1.135670551e-07 wketa=8.233768337e-08 pketa=-1.133313806e-13 dwg=0.0 dwb=0.0 pclm=1.100280049e+00 lpclm=-5.680167483e-07 wpclm=-2.582002469e-06 ppclm=1.609491975e-12 pdiblc1=-2.003109147e-01 lpdiblc1=1.180852641e-06 wpdiblc1=1.886937729e-06 ppdiblc1=-3.774613251e-12 pdiblc2=6.869474325e-03 lpdiblc2=-5.409317078e-09 wpdiblc2=-8.677695359e-09 ppdiblc2=2.630573857e-14 pdiblcb=-4.958541047e-02 lpdiblcb=4.918043384e-08 wpdiblcb=-1.608228360e-09 ppdiblcb=3.217085537e-15 drout=8.601173000e-01 ldrout=-6.003519459e-7 pscbe1=2.355535924e+09 lpscbe1=-3.111680062e+03 wpscbe1=-7.024584736e+03 ppscbe1=1.405191609e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.668768674e-07 lalpha0=-6.738854536e-13 walpha0=-2.037363217e-11 palpha0=4.075523042e-17 alpha1=8.159867060e-01 lalpha1=6.803988720e-8 beta0=1.176738913e+01 lbeta0=4.186039959e-06 wbeta0=-4.702913425e-06 pbeta0=9.407665689e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.611760809e-01 lkt1=9.071521659e-08 wkt1=-9.754508640e-08 pkt1=8.241624584e-14 kt2=-8.754029721e-02 lkt2=6.127258173e-08 wkt2=1.452886480e-07 pkt2=-1.460031677e-13 at=1.573998468e+05 lat=-9.097830411e-02 wat=6.312948634e-02 pat=-8.452587242e-8 ute=-2.580913274e+00 lute=1.591876177e-06 wute=2.599229243e-07 pute=4.510058705e-13 ua1=-8.940665674e-10 lua1=2.875919040e-15 wua1=-2.350730481e-15 pua1=3.896760413e-21 ub1=-3.286796361e-19 lub1=-9.686505929e-25 wub1=4.604046824e-24 pub1=-5.786774035e-30 uc1=1.112783654e-11 luc1=5.766663646e-17 wuc1=4.056478749e-17 puc1=-1.298029296e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.14 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.314468024e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.754687010e-08 wvth0=-1.975606267e-08 pvth0=6.301870618e-14 k1=7.223078201e-01 lk1=-1.083474742e-07 wk1=-2.813131819e-07 pk1=7.146865138e-14 k2=-1.090870399e-01 lk2=4.750147922e-08 wk2=1.606120379e-07 pk2=-6.265970372e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.744605664e+00 ldsub=1.118717944e-06 wdsub=1.291709880e-05 pdsub=-6.794147934e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.067098929e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.097468902e-09 wvoff=-1.896442345e-09 pvoff=-4.533585650e-14 nfactor=2.325140036e+00 lnfactor=3.728254907e-07 wnfactor=9.808660430e-07 pnfactor=-1.200802613e-12 eta0=-4.753090511e-01 leta0=4.830319614e-07 weta0=-6.917910979e-08 peta0=3.461660393e-14 etab=2.469183582e-04 letab=-2.799279117e-10 wetab=-3.866275653e-09 petab=1.934649540e-15 u0=2.824166554e-02 lu0=-2.752296608e-09 wu0=-8.244901712e-09 pu0=7.643537934e-15 ua=-1.263048165e-09 lua=-2.391424758e-16 wua=-8.265299713e-17 pua=5.027183020e-22 ub=2.141316375e-18 lub=8.767931047e-26 wub=-2.550054554e-25 pub=-1.562843116e-31 uc=8.669044640e-11 luc=-4.805367398e-19 wuc=-3.297391807e-16 puc=1.546888282e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.843273509e+05 lvsat=-4.369366421e-02 wvsat=-6.966653454e-01 pvsat=4.179548051e-7 a0=-3.783323516e-01 la0=9.399006038e-07 wa0=8.117649627e-06 pa0=-4.061998814e-12 ags=-1.228154353e+00 lags=1.240046135e-06 wags=1.144234117e-05 pags=-5.725644538e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.234153101e-02 lketa=2.175634589e-08 wketa=-1.450046555e-07 pketa=1.140998492e-13 dwg=0.0 dwb=0.0 pclm=2.513287683e-01 lpclm=2.812664720e-07 wpclm=-3.235909697e-08 ppclm=-9.411483076e-13 pdiblc1=6.615210779e-01 lpdiblc1=3.186836721e-07 wpdiblc1=-1.710014583e-06 ppdiblc1=-1.762545306e-13 pdiblc2=-1.543026337e-03 lpdiblc2=3.006472873e-09 wpdiblc2=4.244205032e-08 ppdiblc2=-2.483399493e-14 pdiblcb=2.417082094e-02 lpdiblcb=-2.460463626e-08 wpdiblcb=3.216456720e-09 ppdiblcb=-1.609485994e-15 drout=1.049590990e+00 ldrout=-7.898997205e-07 wdrout=-7.108420320e-06 pdrout=7.111199712e-12 pscbe1=-1.483910635e+09 lpscbe1=7.292677202e+02 wpscbe1=9.986780585e+03 ppscbe1=-2.966100680e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.128994381e-05 lalpha0=2.099140304e-11 walpha0=1.421457002e-10 palpha0=-1.218276470e-16 alpha1=9.180265880e-01 lalpha1=-3.403989240e-8 beta0=9.611046677e-01 lbeta0=1.499654967e-05 wbeta0=9.331006019e-05 pbeta0=-8.864363100e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.685631945e-01 lkt1=-1.933881430e-09 wkt1=-4.397662358e-10 pkt1=-1.472704250e-14 kt2=-1.712871672e-02 lkt2=-9.166529692e-09 wkt2=3.045405551e-09 pkt2=-3.704308085e-15 at=8.051371031e+04 lat=-1.406210511e-02 wat=-4.977434187e-02 pat=2.842210119e-8 ute=-6.616270746e-01 lute=-3.281604629e-07 wute=2.180573802e-06 pute=-1.470395982e-12 ua1=2.619122030e-09 lua1=-6.386432149e-16 wua1=4.613170050e-15 pua1=-3.069863003e-21 ub1=-1.241180067e-18 lub1=-5.579337394e-26 wub1=-3.422836674e-24 pub1=2.243247975e-30 uc1=1.536964264e-10 luc1=-8.495769773e-17 wuc1=-1.947979223e-16 puc1=1.056518070e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.15 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.137551841e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.363950333e-08 wvth0=1.143094078e-07 pvth0=-4.066448670e-15 k1=2.578512384e-01 lk1=1.240624192e-07 wk1=-3.355262627e-07 pk1=9.859638911e-14 k2=6.454920377e-02 lk2=-3.938453436e-08 wk2=7.623328524e-08 pk2=-2.043733531e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.748036655e-01 ldsub=5.818459021e-08 wdsub=-9.812973617e-07 pdsub=1.604844224e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.014386931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.735129863e-09 wvoff=-1.712052201e-07 pvoff=3.938473212e-14 nfactor=3.036485104e+00 lnfactor=1.687482043e-08 wnfactor=-3.027003159e-06 pnfactor=8.046990646e-13 eta0=0.49 etab=-2.463432642e-04 letab=-3.310423520e-11 wetab=3.539106064e-09 petab=-1.770936822e-15 u0=2.860307686e-02 lu0=-2.933143578e-09 wu0=2.067040832e-08 pu0=-6.825422967e-15 ua=-1.323135195e-09 lua=-2.090754666e-16 wua=1.582794363e-15 pua=-3.306565682e-22 ub=1.932430063e-18 lub=1.922041409e-25 wub=3.095493923e-25 pub=-4.387824764e-31 uc=-3.956346875e-12 luc=4.487830279e-17 wuc=5.865119828e-16 puc=-3.037950078e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.168781891e+04 lvsat=3.768969386e-02 wvsat=3.721284325e-01 pvsat=-1.168599822e-7 a0=1.5 ags=2.482394068e+00 lags=-6.166789003e-07 wags=-4.249483560e-12 pags=2.126403329e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.387472488e-02 lketa=-7.499917695e-09 wketa=6.046346295e-08 pketa=1.128545188e-14 dwg=0.0 dwb=0.0 pclm=1.248389747e+00 lpclm=-2.176538680e-07 wpclm=-4.056794394e-06 ppclm=1.072642895e-12 pdiblc1=3.418493377e+00 lpdiblc1=-1.060880454e-06 wpdiblc1=-1.061063070e-05 ppdiblc1=4.277533667e-12 pdiblc2=6.374537686e-03 lpdiblc2=-9.554049064e-10 wpdiblc2=-1.425354643e-08 ppdiblc2=3.535971429e-15 pdiblcb=6.672051182e-01 lpdiblcb=-3.463732113e-07 wpdiblcb=-3.399586849e-06 ppdiblcb=1.701122663e-12 drout=-2.060339341e+00 ldrout=7.662814279e-07 wdrout=1.421684064e-05 pdrout=-3.559768945e-12 pscbe1=-8.543224250e+08 lpscbe1=4.142274463e+02 wpscbe1=8.124777775e+03 ppscbe1=-2.034371232e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=4.328289667e-05 lalpha0=-1.132026518e-11 walpha0=-2.344130294e-10 palpha0=6.659895226e-17 alpha1=0.85 beta0=4.343426743e+01 lbeta0=-6.256638715e-06 wbeta0=-1.725168945e-04 pbeta0=4.437378467e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.086487723e-01 lkt1=-3.191451909e-08 wkt1=-3.674421612e-07 pkt1=1.689176529e-13 kt2=2.302314085e-03 lkt2=-1.888964263e-08 wkt2=-2.384443201e-07 pkt2=1.171349772e-13 at=8.204118696e+04 lat=-1.482644068e-02 wat=-7.371450278e-03 pat=7.204075861e-9 ute=-1.208490218e+00 lute=-5.451506748e-08 wute=-5.374830147e-06 pute=2.310260156e-12 ua1=1.780566526e-09 lua1=-2.190375874e-16 wua1=-6.885565380e-15 pua1=2.684000718e-21 ub1=-2.179036963e-18 lub1=4.135017759e-25 wub1=3.781134618e-24 pub1=-1.361554424e-30 uc1=-1.484104747e-10 luc1=6.621387661e-17 wuc1=2.124527689e-16 puc1=-9.813277364e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.16 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.765795849e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.433106785e-08 wvth0=4.577582150e-07 pvth0=-9.006293893e-14 k1=4.124772342e-01 lk1=8.534546145e-08 wk1=1.880920012e-07 pk1=-3.251291161e-14 k2=4.255952949e-02 lk2=-3.387851783e-08 wk2=-1.374289433e-07 pk2=3.306176377e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.120434380e+00 ldsub=-1.285146299e-07 wdsub=-1.055935509e-06 pdsub=1.791731426e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.892849404e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.288321112e-08 wvoff=-4.223910930e-07 pvoff=1.022794140e-13 nfactor=3.743685139e+00 lnfactor=-1.602017034e-07 wnfactor=-6.530798722e-06 pnfactor=1.682017940e-12 eta0=1.714692951e+00 leta0=-3.066520927e-07 weta0=-2.888829305e-07 peta0=7.233368585e-14 etab=9.173025369e-02 letab=-2.306321632e-08 wetab=-1.509102451e-07 petab=3.690179067e-14 u0=-2.600543195e-02 lu0=1.074033555e-08 wu0=2.608523595e-08 pu0=-8.181247072e-15 ua=-5.623918542e-09 lua=8.678019763e-16 wua=-1.610170182e-16 pua=1.059781075e-22 ub=4.350834248e-18 lub=-4.133425014e-25 wub=2.891087548e-24 pub=-1.085176397e-30 uc=3.723263434e-10 luc=-4.933949631e-17 wuc=-2.020883903e-15 puc=3.490734555e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.136665712e+05 lvsat=1.465904210e-02 wvsat=2.380270450e-01 pvsat=-8.328220172e-8 a0=1.5 ags=-3.151407387e+00 lags=7.939742800e-07 wags=1.517672701e-11 pags=-2.737744961e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.216582192e-01 lketa=1.698418923e-08 wketa=5.865551833e-07 pketa=-1.204431801e-13 dwg=0.0 dwb=0.0 pclm=1.294324355e+00 lpclm=-2.291554806e-07 wpclm=-3.861756276e-06 ppclm=1.023807106e-12 pdiblc1=-3.890127409e+00 lpdiblc1=7.691324136e-07 wpdiblc1=2.312999512e-05 ppdiblc1=-4.170815371e-12 pdiblc2=-1.066988808e-02 lpdiblc2=3.312365906e-09 wpdiblc2=-2.072601932e-08 ppdiblc2=5.156620387e-15 pdiblcb=-2.464566842e+00 lpdiblcb=4.377943014e-07 wpdiblcb=1.300888967e-05 ppdiblcb=-2.407412181e-12 drout=2.274144656e+00 ldrout=-3.190343545e-07 wdrout=-3.763832674e-06 pdrout=9.424298270e-13 pscbe1=8.212410617e+08 lpscbe1=-5.318570670e+00 wpscbe1=-7.371708867e+01 ppscbe1=1.845809555e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.933005396e-06 lalpha0=-1.467406554e-12 walpha0=3.790852468e-11 palpha0=-1.587913980e-18 alpha1=-3.317959573e+00 lalpha1=1.043619566e-06 walpha1=2.273066027e-05 palpha1=-5.691552755e-12 beta0=4.879438173e+01 lbeta0=-7.598763093e-06 wbeta0=-1.315350603e-04 pbeta0=3.411230222e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-6.211686308e-01 lkt1=7.137674081e-08 wkt1=1.697866138e-06 pkt1=-3.482169574e-13 kt2=-1.670087327e-01 lkt2=2.350431969e-08 wkt2=8.106213789e-07 pkt2=-1.455416322e-13 at=4.052764162e+04 lat=-4.431822545e-03 wat=-2.797783978e-01 pat=7.541232386e-8 ute=-4.588901180e-01 lute=-2.422081862e-07 wute=1.418532112e-05 pute=-2.587425679e-12 ua1=4.757377427e-09 lua1=-9.644042458e-16 wua1=1.311037901e-14 pua1=-2.322803793e-21 ub1=-5.105479826e-18 lub1=1.146256731e-24 wub1=-1.654340121e-26 pub1=-4.106500267e-31 uc1=-1.308406938e-10 luc1=6.181456160e-17 wuc1=7.863898362e-16 puc1=-2.418414499e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.17 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.906260738e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.174171969e-09 wvth0=6.053677575e-07 pvth0=-1.166903719e-13 k1=7.866578881e-01 lk1=1.784663910e-08 wk1=1.371920283e-07 pk1=-2.333101461e-14 k2=3.632657808e-03 lk2=-2.685646052e-08 wk2=-5.593480549e-07 pk2=1.091721742e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.629981589e+00 ldsub=-2.204323606e-07 wdsub=-5.999226392e-06 pdsub=1.070898328e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=7.501412741e-02 lcdscd=-1.255776070e-08 wcdscd=-2.940300821e-07 pcdscd=5.304038054e-14 cit=0.0 voff='6.903011228e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.562335809e-07 wvoff=-3.658396998e-06 pvoff=6.860257552e-13 nfactor=3.549009128e+01 lnfactor=-5.886967654e-06 wnfactor=-1.527429775e-04 pnfactor=2.805737908e-11 eta0=8.400993652e-02 leta0=-1.249155303e-08 weta0=6.798678379e-07 peta0=-1.024202340e-13 etab=4.871470735e-02 letab=-1.530359890e-08 wetab=-3.963140265e-08 petab=1.682808900e-14 u0=7.018040452e-02 lu0=-6.610723675e-09 wu0=1.382630800e-07 pu0=-2.841712055e-14 ua=5.857733218e-09 lua=-1.203384666e-15 wua=8.620350591e-15 pua=-1.478101577e-21 ub=-5.055850015e-18 lub=1.283538679e-24 wub=-2.018586862e-24 pub=-1.995153203e-31 uc=1.867914724e-10 luc=-1.587067540e-17 wuc=4.588799269e-16 puc=-9.825362159e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.218936807e+05 lvsat=-2.290325440e-02 wvsat=-1.602255313e+00 pvsat=2.486881731e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.281788016e+00 lketa=2.262611634e-07 wketa=6.448114199e-06 pketa=-1.177815672e-12 dwg=0.0 dwb=0.0 pclm=-1.025422404e+00 lpclm=1.893059571e-07 wpclm=1.311806618e-05 ppclm=-2.039200047e-12 pdiblc1=-2.196206835e-01 lpdiblc1=1.070060348e-07 wpdiblc1=3.698644863e-06 ppdiblc1=-6.655746675e-13 pdiblc2=-9.575899567e-03 lpdiblc2=3.115020224e-09 wpdiblc2=1.021758303e-07 ppdiblc2=-1.701376716e-14 pdiblcb=-6.671889868e-01 lpdiblcb=1.135635129e-07 wpdiblcb=1.022689933e-06 ppdiblcb=-2.452096241e-13 drout=-3.751154567e-01 ldrout=1.588683264e-07 wdrout=1.379453541e-05 pdrout=-2.224941750e-12 pscbe1=8.187672003e+08 lpscbe1=-4.872308350e+00 wpscbe1=2.767061009e+01 ppscbe1=1.686671823e-7 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.541465026e-05 lalpha0=3.826646397e-12 walpha0=1.750147566e-10 palpha0=-2.632064425e-17 alpha1=1.057523900e+01 lalpha1=-1.462588419e-06 walpha1=-5.303820729e-05 palpha1=7.976469033e-12 beta0=-2.937050130e+01 lbeta0=6.501478322e-06 wbeta0=3.461520388e-04 pbeta0=-5.205815127e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-5.839909174e-01 lkt1=6.467021591e-08 wkt1=7.308639065e-07 pkt1=-1.737784579e-13 kt2=-7.010849465e-02 lkt2=6.024388848e-09 wkt2=1.533319901e-09 pkt2=4.105718345e-16 at=2.529313293e+05 lat=-4.274753616e-02 wat=-1.387331955e+00 pat=2.752050177e-7 ute=-1.083292778e+01 lute=1.629174842e-06 wute=-9.507139222e-07 pute=1.429788175e-13 ua1=-1.561689394e-08 lua1=2.710930941e-15 wua1=1.606143834e-14 pua1=-2.855148337e-21 ub1=9.325143900e-18 lub1=-1.456897914e-24 wub1=-7.659125826e-24 pub1=9.680030595e-31 uc1=2.476838342e-10 luc1=-6.467856515e-18 wuc1=-1.743696895e-15 puc1=2.145634257e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.18 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.164148006e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.470062469e-09 wvth0=-3.884255827e-09 pvth0=3.884271014e-13 k1=5.437797533e-01 lk1=-2.914114662e-07 wk1=-1.619988292e-08 pk1=1.619994626e-12 k2=-2.748715059e-02 lk2=8.768630151e-08 wk2=5.734699003e-09 pk2=-5.734721425e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.061725161e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.039196300e-08 wvoff=2.980634190e-09 pvoff=-2.980645844e-13 nfactor=2.710152389e+00 lnfactor=-2.758249726e-06 wnfactor=2.546847906e-08 pnfactor=-2.546857864e-12 eta0=0.08 etab=-0.07 u0=3.099863670e-02 lu0=1.599639206e-08 wu0=9.286611731e-10 pu0=-9.286648042e-14 ua=-7.591629073e-10 lua=2.436146803e-16 wua=-3.137116100e-17 pua=3.137128366e-21 ub=1.581866692e-18 lub=6.023331977e-25 wub=1.088263642e-25 pub=-1.088267897e-29 uc=5.865943820e-11 luc=-9.417475022e-16 wuc=-4.323207297e-17 puc=4.323224201e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.402701864e+00 la0=-1.894193819e-06 wa0=-1.112945726e-07 pa0=1.112950077e-11 ags=3.729844084e-01 lags=-4.138424618e-07 wags=-2.060712726e-08 pags=2.060720784e-12 a1=0.0 a2=0.42385546 b0=7.668725254e-25 lb0=-7.668755239e-29 wb0=-3.766296555e-30 pb0=3.766311282e-34 b1=2.634188300e-24 lb1=-5.268479596e-29 keta=-9.253996917e-03 lketa=4.593987136e-08 wketa=-9.455522259e-10 pketa=9.455559230e-14 dwg=0.0 dwb=0.0 pclm=1.609390617e-02 lpclm=1.022213380e-06 wpclm=-1.188350296e-08 ppclm=1.188354943e-12 pdiblc1=0.39 pdiblc2=2.777325455e-03 lpdiblc2=2.961344030e-08 wpdiblc2=1.306759243e-09 ppdiblc2=-1.306764352e-13 pdiblcb=-9.299105261e-01 lpdiblcb=9.049140643e-05 wpdiblcb=4.444234582e-06 ppdiblcb=-4.444251959e-10 drout=0.56 pscbe1=8.057324590e+08 lpscbe1=-5.105849865e+03 wpscbe1=-1.769129561e+02 ppscbe1=1.769136478e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.072543108e-01 lkt1=-5.775711810e-07 wkt1=-1.440532921e-08 pkt1=1.440538553e-12 kt2=-4.364567021e-02 lkt2=-1.667673314e-07 wkt2=-7.949455814e-09 pkt2=7.949486896e-13 at=140000.0 ute=-1.761835242e+00 lute=-5.156496004e-06 wute=-1.669302417e-07 pute=1.669308944e-11 ua1=4.313722010e-10 lua1=-5.535241739e-15 wua1=-1.282896440e-16 pua1=1.282901456e-20 ub1=-6.486104031e-19 lub1=8.990438289e-25 wub1=-1.299160521e-25 pub1=1.299165601e-29 uc1=1.485367404e-11 luc1=9.760427809e-17 wuc1=3.323582899e-18 puc1=-3.323595894e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.19 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.163412989e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=1.553671956e-8 k1=5.292094648e-01 wk1=6.479826488e-8 k2=-2.310292122e-02 wk2=-2.293834757e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016530063e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.192230368e-8 nfactor=2.572242599e+00 wnfactor=-1.018719246e-7 eta0=0.08 etab=-0.07 u0=3.179844067e-02 wu0=-3.714572073e-9 ua=-7.469824114e-10 wua=1.254821908e-16 ub=1.611982763e-18 wub=-4.352969467e-25 uc=1.157298363e-11 wuc=1.729249112e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.307994025e+00 wa0=4.451695873e-7 ags=3.522926899e-01 wags=8.242689761e-8 a1=0.0 a2=0.42385546 b0=-3.067430133e-24 wb0=1.506489170e-29 b1=0.0 keta=-6.957048255e-03 wketa=3.782134963e-9 dwg=0.0 dwb=0.0 pclm=6.720357597e-02 wpclm=4.753308259e-8 pdiblc1=0.39 pdiblc2=4.257968523e-03 wpdiblc2=-5.226934785e-9 pdiblcb=3.594571342e+00 wpdiblcb=-1.777659080e-5 drout=0.56 pscbe1=5.504449566e+08 wpscbe1=7.076379900e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.361323053e-01 wkt1=5.762019035e-8 kt2=-5.198387376e-02 wkt2=3.179720162e-8 at=140000.0 ute=-2.019655001e+00 wute=6.677079130e-7 ua1=1.546155246e-10 wua1=5.131485438e-16 ub1=-6.036590905e-19 wub1=5.196540492e-25 uc1=1.973379253e-11 wuc1=-1.329407170e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.20 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.214429505e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.081520778e-08 wvth0=-3.273741878e-08 pvth0=3.862119819e-13 k1=5.145784436e-01 lk1=1.170538901e-07 wk1=9.820608490e-08 pk1=-2.672756226e-13 k2=-1.960026388e-02 lk2=-2.802262825e-08 wk2=-2.196230483e-08 pk2=-7.808723509e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017524766e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.958009487e-10 wvoff=-1.758114517e-08 pvoff=4.527294454e-14 nfactor=2.037542839e+00 lnfactor=4.277807153e-06 wnfactor=1.676306533e-06 pnfactor=-1.422612293e-11 eta0=0.08 etab=-0.07 u0=3.296822585e-02 lu0=-9.358738773e-09 wu0=-7.690467856e-09 pu0=3.180872084e-14 ua=-6.533344060e-10 lua=-7.492206594e-16 wua=-2.967403534e-16 pua=3.377945443e-21 ub=1.572654670e-18 lub=3.146401164e-25 wub=-1.532449980e-25 pub=-2.256525872e-30 uc=-1.013326580e-10 luc=9.032892790e-16 wuc=5.316849805e-16 puc=-2.870220829e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.064900943e+00 la0=1.944839705e-06 wa0=1.510896977e-06 pa0=-8.526235817e-12 ags=2.099268989e-01 lags=1.138981992e-06 wags=4.961602859e-07 pags=-3.310028876e-12 a1=0.0 a2=0.42385546 b0=-6.135160108e-24 lb0=2.454303928e-29 wb0=3.013125600e-29 pb0=-1.205368053e-34 b1=0.0 keta=-9.999992786e-03 lketa=2.434474604e-08 wketa=-1.833946167e-09 pketa=4.493084493e-14 dwg=0.0 dwb=0.0 pclm=-3.579713867e-01 lpclm=3.401565945e-06 wpclm=1.052232518e-07 ppclm=-4.615439103e-13 pdiblc1=0.39 pdiblc2=5.657438365e-03 lpdiblc2=-1.119630593e-08 wpdiblc2=-1.229612468e-08 ppdiblc2=5.655628318e-14 pdiblcb=7.214496497e+00 lpdiblcb=-2.896081663e-05 wpdiblcb=-3.555491925e-05 ppdiblcb=1.422335790e-10 drout=0.56 pscbe1=3.034901470e+08 lpscbe1=1.975735036e+03 wpscbe1=1.407704225e+03 ppscbe1=-5.600803605e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.571936509e-01 lkt1=1.684990000e-07 wkt1=1.253984533e-07 pkt1=-5.422526049e-13 kt2=-6.235832228e-02 lkt2=8.299964454e-08 wkt2=6.520270516e-08 pkt2=-2.672570899e-13 at=140000.0 ute=-2.360816710e+00 lute=2.729427067e-06 wute=1.581427534e-06 pute=-7.310114231e-12 ua1=-4.808083547e-10 lua1=5.083639485e-15 wua1=2.491844488e-15 pua1=-1.583034123e-20 ub1=-1.855114199e-19 lub1=-3.345344861e-24 wub1=-9.143566132e-25 pub1=1.147264600e-29 uc1=2.758544161e-11 luc1=-6.281626264e-17 wuc1=-7.104339671e-17 puc1=4.620171801e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.21 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.902585930e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.393441518e-08 wvth0=1.273673423e-07 pvth0=-2.542696632e-13 k1=5.392881432e-01 lk1=1.820543048e-08 wk1=2.345025689e-09 pk1=1.162060959e-13 k2=-1.986551524e-02 lk2=-2.696151910e-08 wk2=-2.871039032e-08 pk2=1.918625693e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.296830322e+00 ldsub=-2.947609389e-06 wdsub=-2.145091381e-06 pdsub=8.581204254e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.066154553e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.024961738e-08 wvoff=3.789037041e-10 pvoff=-2.657427333e-14 nfactor=3.451899107e+00 lnfactor=-1.380170934e-06 wnfactor=-3.872666475e-06 pnfactor=7.971938752e-12 eta0=2.752600354e-01 leta0=-7.811164882e-07 weta0=-5.684492159e-07 peta0=2.274019127e-12 etab=-2.406990244e-01 letab=6.828628408e-07 wetab=4.969461691e-07 petab=-1.987978982e-12 u0=3.136212758e-02 lu0=-2.933717721e-09 wu0=5.000156996e-09 pu0=-1.895874060e-14 ua=-8.528743887e-10 lua=4.901729144e-17 wua=9.911510278e-16 pua=-1.774123648e-21 ub=1.713934631e-18 lub=-2.505349677e-25 wub=-8.558227277e-25 pub=5.540597547e-31 uc=1.658611426e-10 luc=-1.655903961e-16 wuc=-3.163932560e-16 puc=5.224237150e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.296171895e+00 la0=-2.980725529e-06 wa0=-3.509334004e-06 pa0=1.155665102e-11 ags=5.459549050e-01 lags=-2.052614186e-07 wags=-1.121424763e-06 pags=3.160943795e-12 a1=0.0 a2=0.42385546 b0=3.068029816e-24 lb0=-1.227331886e-29 wb0=-1.506783689e-29 pb0=6.027723908e-35 b1=0.0 keta=-1.066714159e-02 lketa=2.701360211e-08 wketa=2.592489432e-08 pketa=-6.611537072e-14 dwg=0.0 dwb=0.0 pclm=6.025325291e-01 lpclm=-4.408252756e-07 wpclm=-3.752460009e-07 ppclm=1.460520964e-12 pdiblc1=0.39 pdiblc2=3.101284362e-04 lpdiblc2=1.019502459e-08 wpdiblc2=5.307527020e-09 ppdiblc2=-1.386520663e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.826104865e+08 lpscbe1=5.906634211e+01 wpscbe1=7.490559788e+01 ppscbe1=-2.690879728e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.953020551e-01 lkt1=-7.909158272e-08 wkt1=-5.734345830e-08 pkt1=1.887864936e-13 kt2=-4.019663021e-02 lkt2=-5.655788958e-09 wkt2=-7.314905443e-09 pkt2=2.284170692e-14 at=1.622768398e+05 lat=-8.911606945e-02 wat=7.650825925e-03 pat=-3.060629517e-8 ute=-1.524142064e+00 lute=-6.175986579e-07 wute=-1.211928552e-06 pute=3.864402316e-12 ua1=1.242815922e-09 lua1=-1.811531558e-15 wua1=-3.541988009e-15 pua1=8.307347992e-21 ub1=-1.496596327e-18 lub1=1.899507400e-24 wub1=3.501937242e-24 pub1=-6.194256193e-30 uc1=3.120698193e-12 luc1=3.505227676e-17 wuc1=1.837167575e-17 puc1=1.043219289e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.22 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.332224896e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.010176900e-09 wvth0=-1.300652481e-07 pvth0=2.606961737e-13 k1=4.312570044e-01 lk1=2.343099483e-07 wk1=5.837452191e-07 pk1=-1.046821618e-12 k2=4.357746534e-03 lk2=-7.541751395e-08 wk2=-1.825731576e-07 pk2=3.269719519e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.500214865e+00 ldsub=2.647574630e-06 wdsub=6.871498134e-06 pdsub=-9.455500262e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.463644626e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.371699452e-08 wvoff=4.824463636e-08 pvoff=-1.223244541e-13 nfactor=2.507695437e+00 lnfactor=5.086055905e-07 wnfactor=2.008417883e-06 pnfactor=-3.792529468e-12 eta0=-2.280162057e-01 leta0=2.256327751e-07 weta0=1.122328176e-06 peta0=-1.108196750e-12 etab=7.955202580e-02 letab=4.223552229e-08 wetab=-3.935166719e-07 petab=-2.067051293e-13 u0=3.282442487e-02 lu0=-5.858884067e-09 wu0=-1.093246478e-09 pu0=-6.769551130e-15 ua=-3.285700639e-10 lua=-9.997963611e-16 wua=6.440202226e-16 pua=-1.079726309e-21 ub=1.013225334e-18 lub=1.151157603e-24 wub=-1.066025960e-24 pub=9.745484090e-31 uc=1.510350620e-10 luc=-1.359324379e-16 wuc=-2.844087529e-16 puc=4.584422028e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.406886462e+04 lvsat=3.186849984e-02 wvsat=5.923754944e-02 pvsat=-1.184982608e-7 a0=-4.075307497e-01 la0=2.427736907e-06 wa0=7.641453719e-06 pa0=-1.074928439e-11 ags=-3.349586523e-01 lags=1.556910133e-06 wags=1.141096424e-06 pags=-1.364983225e-12 a1=0.0 a2=0.42385546 b0=-6.136059632e-24 lb0=6.138458831e-30 wb0=3.013567378e-29 pb0=-3.014745683e-35 b1=0.0 keta=9.528481514e-02 lketa=-1.849317386e-07 wketa=-1.256820769e-07 pketa=2.371578501e-13 dwg=0.0 dwb=0.0 pclm=1.238015435e+00 lpclm=-1.712039561e-06 wpclm=-3.258454284e-06 ppclm=7.228064864e-12 pdiblc1=2.196427337e-01 lpdiblc1=3.407811422e-07 wpdiblc1=-1.755562671e-07 ppdiblc1=3.511811766e-13 pdiblc2=3.187179521e-03 lpdiblc2=4.439797488e-09 wpdiblc2=9.406945540e-09 ppdiblc2=-2.206564654e-14 pdiblcb=-5.005092380e-02 lpdiblcb=5.011164250e-08 wpdiblcb=6.780202251e-10 ppdiblcb=-1.356305556e-15 drout=8.601173000e-01 ldrout=-6.003519459e-7 pscbe1=5.780143354e+08 lpscbe1=4.683386413e+02 wpscbe1=1.705253944e+03 ppscbe1=-3.530422131e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-9.287635897e-06 lalpha0=1.863891499e-11 walpha0=2.704201641e-11 palpha0=-5.409460625e-17 alpha1=1.088294264e+00 lalpha1=-4.766817003e-07 walpha1=-1.337368314e-06 palpha1=2.675259539e-12 beta0=7.344075289e+00 lbeta0=1.303439715e-05 wbeta0=1.702105127e-05 pbeta0=-3.404875777e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.689871834e-01 lkt1=6.830748474e-08 wkt1=-5.918287173e-08 pkt1=1.924660396e-13 kt2=-7.332560461e-02 lkt2=6.061511328e-08 wkt2=7.547685272e-08 pkt2=-1.427741810e-13 at=1.784994087e+05 lat=-1.215675504e-01 wat=-4.049556828e-02 pat=6.570531849e-8 ute=-3.299654754e+00 lute=2.934120948e-06 wute=3.789836271e-06 pute=-6.141083022e-12 ua1=-2.584024079e-09 lua1=5.843644738e-15 wua1=5.949059827e-15 pua1=-1.067845868e-20 ub1=5.721107566e-19 lub1=-2.238715630e-24 wub1=1.800472146e-25 pub1=4.508227203e-31 uc1=-1.051621193e-10 luc1=2.516602503e-16 wuc1=6.116929027e-16 puc1=-1.082552514e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.23 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.631332819e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.810643573e-08 wvth0=3.157481685e-07 pvth0=-1.852915560e-13 k1=9.986117363e-01 lk1=-3.332666194e-07 wk1=-1.638308580e-06 pk1=1.176101004e-12 k2=-1.860580729e-01 lk2=1.150727580e-07 wk2=5.386354079e-07 pk2=-3.945186062e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.897783229e+00 ldsub=-7.517520810e-07 wdsub=-4.971554508e-06 pdsub=2.392183014e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-7.649949018e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.185713214e-08 wvoff=-1.502670412e-07 pvoff=7.626484151e-14 nfactor=3.380303252e+00 lnfactor=-3.643434140e-07 wnfactor=-4.201295860e-06 pnfactor=2.419612273e-12 eta0=-4.953283500e-01 leta0=4.930494384e-07 weta0=2.914051193e-08 peta0=-1.458164990e-14 etab=2.434948130e-01 letab=-1.217713665e-07 wetab=-1.198515552e-06 petab=5.986085054e-13 u0=2.703631762e-02 lu0=-6.851366283e-11 wu0=-2.325146351e-09 pu0=-5.537169584e-15 ua=-1.161794829e-09 lua=-1.662458056e-16 wua=-5.799326347e-16 pua=1.447051136e-22 ub=2.017074445e-18 lub=1.469159879e-25 wub=3.551767282e-25 pub=-4.472099695e-31 uc=-5.962263353e-11 luc=7.480762478e-17 wuc=3.888397626e-16 puc=-2.150695528e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.848607431e+04 lvsat=1.744565302e-02 wvsat=-1.768532223e-01 pvsat=1.176848225e-7 a0=2.538920626e+00 la0=-5.198665308e-07 wa0=-6.209685720e-06 pa0=3.107270847e-12 ags=1.097100114e+00 lags=1.242914316e-07 wags=2.245376730e-08 pags=-2.459031790e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.770671126e-01 lketa=8.752667874e-08 wketa=3.202155991e-07 pketa=-2.089141719e-13 dwg=0.0 dwb=0.0 pclm=-1.406054435e+00 lpclm=9.330641403e-07 wpclm=8.107450903e-06 ppclm=-4.142284392e-12 pdiblc1=-3.095184037e-01 lpdiblc1=8.701491817e-07 wpdiblc1=3.058995303e-06 ppdiblc1=-2.884635103e-12 pdiblc2=9.472470713e-03 lpdiblc2=-1.847951252e-09 wpdiblc2=-1.165772144e-08 ppdiblc2=-9.927432770e-16 pdiblcb=2.510184759e-02 lpdiblcb=-2.507051362e-08 wpdiblcb=-1.356040450e-09 ppdiblcb=6.785504369e-16 drout=-2.772720638e-01 ldrout=5.374821372e-07 wdrout=-5.918747599e-07 pdrout=5.921061829e-13 pscbe1=1.292532361e+09 lpscbe1=-2.464587605e+02 wpscbe1=-3.649002865e+03 ppscbe1=1.825928193e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.334146913e-05 lalpha0=-1.400294802e-11 walpha0=-7.704996959e-11 palpha0=5.003807972e-17 alpha1=3.734114727e-01 lalpha1=2.384806098e-07 walpha1=2.674736628e-06 palpha1=-1.338414136e-12 beta0=3.294905457e+01 lbeta0=-1.258059368e-05 wbeta0=-6.379050288e-05 pbeta0=4.679439370e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.239013681e-01 lkt1=2.320404084e-08 wkt1=2.713393958e-07 pkt1=-1.381854621e-13 kt2=1.002820824e-02 lkt2=-2.277129092e-08 wkt2=-1.303288249e-07 pkt2=6.311196666e-14 at=4.956000564e+04 lat=7.422268057e-03 wat=1.022467926e-01 pat=-7.709285464e-8 ute=1.057862942e+00 lute=-1.425100538e-06 wute=-6.264257788e-06 pute=3.916942188e-12 ua1=5.496093080e-09 lua1=-2.239631747e-15 wua1=-9.516331001e-15 pua1=4.792979116e-21 ub1=-1.382578441e-18 lub1=-2.832621492e-25 wub1=-2.728395042e-24 pub1=3.360402178e-30 uc1=4.000687126e-10 luc1=-2.537681269e-16 wuc1=-1.404791842e-15 puc1=9.347206766e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.24 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.617437358e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.127644791e-08 wvth0=-1.213739826e-07 pvth0=3.344043431e-14 k1=-8.066555269e-02 lk1=2.067940226e-07 wk1=1.327011619e-06 pk1=-3.077185362e-13 k2=1.770284158e-01 lk2=-6.661245312e-08 wk2=-4.761793450e-07 pk2=1.132855629e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.047128088e-01 ldsub=4.540601954e-08 wdsub=-6.370642028e-07 pdsub=2.232430754e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.399405904e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.117765790e-10 wvoff=1.788691482e-08 pvoff=-7.877884708e-15 nfactor=2.217924014e+00 lnfactor=2.173006950e-07 wnfactor=9.931484474e-07 pnfactor=-1.796409086e-13 eta0=0.49 etab=2.074390464e-03 letab=-9.667598663e-10 wetab=-7.858578894e-09 petab=2.814471927e-15 u0=3.696083797e-02 lu0=-5.034654326e-09 wu0=-2.037657905e-08 pu0=3.495604878e-15 ua=-8.475116429e-10 lua=-3.235102831e-16 wua=-7.531080024e-16 pua=2.313605090e-22 ub=2.038900016e-18 lub=1.359946685e-25 wub=-2.133503136e-25 pub=-1.627241545e-31 uc=1.711665017e-10 luc=-4.067718138e-17 wuc=-2.735587062e-16 puc=1.163886794e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.055039093e+05 lvsat=3.926171526e-03 wvsat=-3.951267109e-02 pvsat=4.896084673e-8 a0=1.5 ags=2.673519658e+00 lags=-6.645347204e-07 wags=-9.386682737e-07 pags=2.350336402e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.703407186e-02 lketa=-9.599807032e-09 wketa=-1.404495377e-07 pketa=2.159851659e-14 dwg=0.0 dwb=0.0 pclm=3.402336774e-01 lpclm=5.923728531e-08 wpclm=4.033798356e-07 ppclm=-2.872365662e-13 pdiblc1=1.859010953e+00 lpdiblc1=-2.149633914e-07 wpdiblc1=-2.951635112e-06 ppdiblc1=1.230302610e-13 pdiblc2=9.103916561e-03 lpdiblc2=-1.663530072e-09 wpdiblc2=-2.765818660e-08 ppdiblc2=7.013745484e-15 pdiblcb=-3.165795182e-01 lpdiblcb=1.459037667e-07 wpdiblcb=1.432017576e-06 ppdiblcb=-7.165687071e-13 drout=5.933867677e-01 ldrout=1.018122939e-07 wdrout=1.183749520e-06 pdrout=-2.964002260e-13 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.554886287e-05 lalpha0=5.457424100e-12 walpha0=5.452397900e-11 palpha0=-1.580033999e-17 alpha1=0.85 beta0=-4.210918751e+00 lbeta0=6.013922529e-06 wbeta0=6.148014503e-05 pbeta0=-1.588991108e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.417881835e-01 lkt1=-1.788465768e-08 wkt1=-2.046864928e-07 pkt1=1.000136083e-13 kt2=-3.094003958e-02 lkt2=-2.271148424e-09 wkt2=-7.518307660e-08 pkt2=3.551753052e-14 at=9.510846684e+04 lat=-1.536977200e-02 wat=-7.154802405e-02 pat=9.872507447e-9 ute=-2.413220214e+00 lute=3.117982335e-07 wute=5.418904064e-07 pute=5.112068872e-13 ua1=1.376616976e-09 lua1=-1.782829795e-16 wua1=-4.901671383e-15 pua1=2.483844976e-21 ub1=-3.878633954e-18 lub1=9.657415651e-25 wub1=1.212826674e-23 pub1=-4.073737670e-30 uc1=-3.358003181e-10 luc1=1.144541133e-16 wuc1=1.132769639e-15 puc1=-3.350522502e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.25 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='7.756382543e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.979461029e-08 wvth0=-5.198670828e-07 pvth0=1.332195202e-13 k1=4.539393353e-01 lk1=7.293377005e-08 wk1=-1.553841127e-08 pk1=2.844390850e-14 k2=-8.673340762e-03 lk2=-2.011440459e-08 wk2=1.141880808e-07 pk2=-3.453712727e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=9.578166023e-01 ldsub=-1.181252924e-07 wdsub=-2.572802510e-07 pdsub=1.281485919e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-7.158870662e-03 lcdscd=3.144628184e-09 wcdscd=6.167965307e-08 pcdscd=-1.544403001e-14 cit=0.0 voff='-2.589623018e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.969018876e-08 wvoff=6.091357650e-07 pvoff=-1.559212756e-13 nfactor=-1.018394649e+00 lnfactor=1.027645761e-06 wnfactor=1.685692754e-05 pnfactor=-4.151788419e-12 eta0=1.517477597e+00 leta0=-2.572711429e-07 weta0=6.796894011e-07 peta0=-1.701881088e-13 etab=-3.885904740e-02 letab=9.282604575e-09 wetab=4.904454151e-07 petab=-1.219563634e-13 u0=-2.246823902e-02 lu0=9.845851689e-09 wu0=8.713225448e-09 pu0=-3.788220361e-15 ua=-7.469116758e-09 lua=1.334480043e-15 wua=8.901197961e-15 pua=-2.185990816e-21 ub=7.816025157e-18 lub=-1.310545473e-24 wub=-1.412730358e-23 pub=3.321204518e-30 uc=-2.595059472e-10 luc=6.715932377e-17 wuc=1.082197380e-15 puc=-2.230804427e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.350635952e+05 lvsat=-3.475307767e-03 wvsat=1.329410823e-01 pvsat=5.779978974e-9 a0=1.5 ags=-3.151402995e+00 lags=7.939734877e-07 wags=-6.392935609e-12 pags=1.153228047e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.205248154e-02 lketa=-8.352461652e-09 wketa=-7.013042587e-08 pketa=3.991243853e-15 dwg=0.0 dwb=0.0 pclm=5.321809301e-01 lpclm=1.117542075e-08 wpclm=-1.186854768e-07 ppclm=-1.565161106e-13 pdiblc1=2.542229155e+00 lpdiblc1=-3.860350803e-07 wpdiblc1=-8.460864600e-06 ppdiblc1=1.502491742e-12 pdiblc2=-1.847253556e-02 lpdiblc2=5.241365350e-09 wpdiblc2=1.759467069e-08 ppdiblc2=-4.317162705e-15 pdiblcb=1.236449033e+00 lpdiblcb=-2.429606053e-07 wpdiblcb=-5.167694939e-06 ppdiblcb=9.359399094e-13 drout=3.838008024e-01 ldrout=1.542907333e-07 wdrout=5.520103454e-06 pdrout=-1.382184224e-12 pscbe1=7.831160832e+08 lpscbe1=4.227580821e+00 wpscbe1=1.135239070e+02 ppscbe1=-2.842536459e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.154240320e-05 lalpha0=-1.325985103e-12 walpha0=5.369305880e-13 palpha0=-2.282468951e-18 alpha1=1.980401078e+00 lalpha1=-2.830422563e-07 walpha1=-3.290871095e-06 palpha1=8.240045044e-13 beta0=7.916927103e+00 lbeta0=2.977219078e-06 wbeta0=6.922401175e-05 pbeta0=-1.782890561e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.352730142e-01 lkt1=5.523102551e-09 wkt1=2.937635779e-07 pkt1=-2.479380334e-14 kt2=-2.403456685e-02 lkt2=-4.000216647e-09 wkt2=1.084406506e-07 pkt2=-1.046019816e-14 at=1.255163911e+05 lat=-2.298364257e-02 wat=-6.971787140e-01 pat=1.665248015e-7 ute=2.478595444e+00 lute=-9.130683810e-07 wute=-2.413813483e-07 pute=7.073310851e-13 ua1=5.712557732e-09 lua1=-1.263963521e-15 wua1=8.419257377e-15 pua1=-8.515956977e-22 ub1=-2.370881291e-18 lub1=5.882138680e-25 wub1=-1.344681858e-23 pub1=2.330033519e-30 uc1=3.596936738e-10 luc1=-5.969132282e-17 wuc1=-1.622743152e-15 puc1=3.549033530e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.26 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.140268049e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.260225932e-08 wvth0=4.904411039e-07 pvth0=-4.903098395e-14 k1=6.799744235e-01 lk1=3.215907445e-08 wk1=6.611403405e-07 pk1=-9.362284821e-14 k2=-8.974239384e-02 lk2=-5.490277036e-09 wk2=-1.007605795e-07 pk2=4.237676513e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.353763174e-01 ldsub=-5.842666978e-09 wdsub=3.588933925e-07 pdsub=1.699641219e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=3.420427281e-02 lcdscd=-4.316910629e-09 wcdscd=-9.360304699e-08 pcdscd=1.256757153e-14 cit=0.0 voff='1.309006814e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.063758463e-08 wvoff=-9.110460551e-07 pvoff=1.183058432e-13 nfactor=1.179678852e+01 lnfactor=-1.284097945e-06 wnfactor=-3.637943381e-05 pnfactor=5.451572041e-12 eta0=5.452200696e-01 leta0=-8.188463534e-08 weta0=-1.585246739e-06 peta0=2.383859863e-13 etab=1.742801830e-01 letab=-2.916579435e-08 wetab=-6.563138406e-07 petab=8.490868546e-14 u0=2.030045638e-01 lu0=-3.082741268e-08 wu0=-5.140685096e-07 pu0=9.051689961e-14 ua=2.038261358e-08 lua=-3.689721444e-15 wua=-6.271485190e-14 pua=1.073290003e-20 ub=-1.645359317e-17 lub=3.067475247e-24 wub=5.395848804e-23 pub=-8.960859519e-30 uc=6.011716828e-10 luc=-8.809917459e-17 wuc=-1.576241566e-15 puc=2.564780172e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.695953836e+05 lvsat=5.148243007e-02 wvsat=8.115664221e-01 pvsat=-1.166379247e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.549722093e-01 lketa=-1.243293943e-07 wketa=-3.063783964e-06 pketa=5.440193993e-13 dwg=0.0 dwb=0.0 pclm=2.970625506e+00 lpclm=-4.286980348e-07 wpclm=-6.507492153e-06 ppclm=9.959671145e-13 pdiblc1=7.904011109e-01 lpdiblc1=-7.002106763e-08 wpdiblc1=-1.261816595e-06 ppdiblc1=2.038482730e-13 pdiblc2=1.533702176e-02 lpdiblc2=-8.575745043e-10 wpdiblc2=-2.017755531e-08 ppdiblc2=2.496606915e-15 pdiblcb=-9.766588286e-01 lpdiblcb=1.562641350e-07 wpdiblcb=2.542571217e-06 ppdiblcb=-4.549227128e-13 drout=5.243473457e+00 ldrout=-7.223504765e-07 wdrout=-1.379971444e-05 pdrout=2.102937046e-12 pscbe1=8.724098391e+08 lpscbe1=-1.188020911e+01 wpscbe1=-2.357813706e+02 ppscbe1=3.458616374e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.505496078e-05 lalpha0=-3.763528876e-12 walpha0=-7.285371686e-11 palpha0=1.095654333e-17 alpha1=-1.787602515e+00 lalpha1=3.966716799e-07 walpha1=7.678699222e-06 palpha1=-1.154807255e-12 beta0=7.736474050e+01 lbeta0=-9.550541429e-06 wbeta0=-1.780505636e-04 pbeta0=2.677720231e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-7.033246839e-01 lkt1=7.191631131e-08 wkt1=1.316940913e-06 pkt1=-2.093657860e-13 kt2=-1.293564417e-01 lkt2=1.499890168e-08 wkt2=2.925143260e-07 pkt2=-4.366543254e-14 at=-2.922389739e+05 lat=5.237566549e-02 wat=1.290131335e+00 pat=-1.919680455e-7 ute=-2.515689494e+01 lute=4.072125364e-06 wute=6.939775516e-05 pute=-1.185494239e-11 ua1=-3.028374087e-08 lua1=5.229444780e-15 wua1=8.809387298e-14 pua1=-1.522417928e-20 ub1=1.803923590e-17 lub1=-3.093587582e-24 wub1=-5.045614044e-23 pub1=9.006182099e-30 uc1=-4.778782195e-10 luc1=9.139910857e-17 wuc1=1.819713936e-15 puc1=-2.660849236e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.27 nmos lmin=2.0e-05 lmax=0.0001 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.076632539e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.803024017e-07 wvth0=2.159361438e-08 pvth0=-4.318807307e-13 k1=5.345415456e-01 lk1=3.385239066e-07 wk1=1.069477533e-08 pk1=-2.138996882e-13 k2=-2.273832376e-02 lk2=-1.648797882e-07 wk2=-8.090285111e-09 pk2=1.618088655e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.079869812e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.477509904e-08 wvoff=8.262981167e-09 pvoff=-1.652628542e-13 nfactor=3.032035046e+00 lnfactor=-9.895894376e-06 wnfactor=-9.116098292e-07 pnfactor=1.823255302e-11 eta0=0.08 etab=-0.07 u0=3.159595381e-02 lu0=-2.146949599e-08 wu0=-8.102734806e-10 pu0=1.620578643e-14 ua=-8.542591606e-10 lua=3.007646410e-15 wua=2.454770457e-16 pua=-4.909636895e-21 ub=1.773438164e-18 lub=-6.219684878e-24 wub=-4.488845531e-25 pub=8.977866576e-30 uc=4.968409686e-11 luc=4.257663863e-16 wuc=-1.710268231e-17 puc=3.420603333e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.328930550e+00 la0=2.639600605e-06 wa0=1.034715757e-07 pa0=-2.069471972e-12 ags=3.653564583e-01 lags=3.049967966e-07 wags=1.599681550e-09 pags=-3.199425647e-14 a1=0.0 a2=0.42385546 b0=-5.268352994e-25 lb0=5.268373594e-29 b1=7.668759614e-24 lb1=-1.533781908e-28 wb1=-1.465685546e-29 pb1=2.931428401e-34 keta=-1.580862553e-02 lketa=2.030184795e-07 wketa=1.813655788e-08 pketa=-3.627382491e-13 dwg=0.0 dwb=0.0 pclm=-1.087933307e-01 lpclm=3.846561813e-06 wpclm=3.516934663e-07 ppclm=-7.034006838e-12 pdiblc1=0.39 pdiblc2=2.938954653e-03 lpdiblc2=-9.528533337e-09 wpdiblc2=8.362175333e-10 ppdiblc2=-1.672467763e-14 pdiblcb=5.966663033e-01 lpdiblcb=-6.216687341e-05 wpdiblcb=2.220446049e-22 ppdiblcb=-6.661338148e-27 drout=0.56 pscbe1=8.886509661e+08 lpscbe1=-1.902740919e+03 wpscbe1=-4.183087964e+02 ppscbe1=8.366339487e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.850388507e-01 lkt1=-6.260352250e-07 wkt1=-7.907990965e-08 pkt1=1.581629113e-12 kt2=-4.590762382e-02 lkt2=9.692113127e-08 wkt2=-1.364361439e-09 pkt2=2.728776224e-14 at=140000.0 ute=-1.651224065e+00 lute=-2.781573069e-06 wute=-4.889461432e-07 pute=9.779114043e-12 ua1=6.666343311e-10 lua1=-6.715217902e-15 wua1=-8.131946382e-16 pua1=1.626421072e-20 ub1=-1.031933345e-18 lub1=1.213570416e-23 wub1=9.860297970e-25 pub1=-1.972098148e-29 uc1=1.313509320e-11 luc1=4.064557052e-17 wuc1=8.326787595e-18 puc1=-1.665390077e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.28 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.5216781+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.030982152 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.53725 eta0=0.08 etab=-0.07 u0=0.0305225 ua=-7.0387978e-10 ub=1.46246e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.460908 ags=0.380606 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.29 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.101977779e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.184706554e-8 k1=5.483118416e-01 lk1=2.524578124e-8 k2=-2.714422788e-02 lk2=-3.070489359e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077915297e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.634687659e-8 nfactor=2.613347438e+00 lnfactor=-6.088092565e-7 eta0=0.08 etab=-0.07 u0=3.032658085e-02 lu0=1.567429798e-9 ua=-7.552635323e-10 lua=4.110901092e-16 ub=1.520015626e-18 lub=-4.604675083e-25 uc=8.129900937e-11 luc=-8.262011279e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.583888020e+00 la0=-9.838882462e-7 ags=3.803559756e-01 lags=2.000293260e-9 a1=0.0 a2=0.42385546 b0=4.214805989e-24 lb0=-1.686087194e-29 b1=0.0 keta=-1.062994597e-02 lketa=3.977831183e-8 dwg=0.0 dwb=0.0 pclm=-3.218276199e-01 lpclm=3.243027455e-06 wpclm=-1.110223025e-22 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=1.433768648e-03 lpdiblc2=8.230551467e-9 pdiblcb=-4.998476267e+00 lpdiblcb=1.989584970e-5 drout=0.56 pscbe1=7.870309262e+08 lpscbe1=5.188136624e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141197830e-01 lkt1=-1.776260414e-8 kt2=-3.996145347e-02 lkt2=-8.802098461e-9 at=140000.0 ute=-1.817602669e+00 lute=2.184320239e-7 ua1=3.751302750e-10 lua1=-3.540195022e-16 wua1=4.135903063e-31 ub1=-4.995892647e-19 lub1=5.954632198e-25 uc1=3.182318579e-12 luc1=9.588479350e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.30 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.340087664e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.406198640e-9 k1=5.400936501e-01 lk1=5.812176032e-8 k2=-2.972741965e-02 lk2=-2.037111647e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064853034e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.112146062e-8 nfactor=2.121653639e+00 lnfactor=1.358158189e-6 eta0=0.08 etab=-0.07 u0=3.307966154e-02 lu0=-9.445969399e-9 ua=-5.124179691e-10 lua=-5.603870960e-16 ub=1.419962942e-18 lub=-6.021765480e-26 uc=5.718132279e-11 luc=1.386006354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.090729680e+00 la0=9.889379399e-7 ags=1.607499777e-01 lags=8.805101507e-7 a1=0.0 a2=0.42385546 b0=-2.107711977e-24 lb0=8.431672024e-30 b1=0.0 keta=-1.762043929e-03 lketa=4.303236316e-09 pketa=1.734723476e-30 dwg=0.0 dwb=0.0 pclm=4.736370264e-01 lpclm=6.085784249e-8 pdiblc1=0.39 pdiblc2=2.133242770e-03 lpdiblc2=5.432381483e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.083402602e+08 lpscbe1=-3.336430185e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.149993040e-01 lkt1=-1.424417615e-8 kt2=-4.270927102e-02 lkt2=2.190246143e-9 at=1.649048679e+05 lat=-9.962920960e-2 ute=-1.940434682e+00 lute=7.098081038e-7 ua1=2.615718673e-11 lua1=1.042009300e-15 ub1=-2.936948702e-19 lub1=-2.281948629e-25 uc1=9.431295441e-12 luc1=7.088644271e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.31 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.885455964e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.753791758e-8 k1=6.317711558e-01 lk1=-1.252690968e-7 k2=-5.835540395e-02 lk2=3.689604566e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.806460635e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.573495597e-8 nfactor=3.197578958e+00 lnfactor=-7.941131350e-7 eta0=1.574990403e-01 leta0=-1.550283827e-7 etab=-5.561937937e-02 letab=-2.876686407e-8 u0=3.244889907e-02 lu0=-8.184197843e-9 ua=-1.073516895e-10 lua=-1.370678036e-15 ub=6.470496747e-19 lub=1.485911089e-24 uc=5.334179128e-11 luc=2.154062782e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.441672627e+04 lvsat=-8.835179470e-3 a0=2.217278084e+00 la0=-1.264599349e-6 ags=5.700341213e-02 lags=1.088043847e-6 a1=0.0 a2=0.42385546 b0=4.215423954e-24 lb0=-4.217072185e-30 b1=0.0 keta=5.211352366e-02 lketa=-1.034689642e-07 wketa=2.515349040e-23 pketa=9.540979118e-30 dwg=0.0 dwb=0.0 pclm=1.187494024e-01 lpclm=7.707718516e-7 pdiblc1=1.593398571e-01 lpdiblc1=4.614104738e-7 pdiblc2=6.418427744e-03 lpdiblc2=-3.139663973e-9 pdiblcb=-4.981802656e-02 lpdiblcb=4.964575696e-8 drout=8.601173000e-01 ldrout=-6.003519459e-7 pscbe1=1.163762255e+09 lpscbe1=-7.443472606e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.188739200e-09 lalpha0=5.763378680e-14 alpha1=6.289135890e-01 lalpha1=4.422592668e-7 beta0=1.319073842e+01 lbeta0=1.338784839e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.893162635e-01 lkt1=1.344188007e-07 wkt1=4.440892099e-22 kt2=-4.739960715e-02 lkt2=1.157275232e-08 wkt2=-5.551115123e-23 at=1.645893428e+05 lat=-9.899803587e-2 ute=-1.997861131e+00 lute=8.246834563e-7 ua1=-5.405457877e-10 lua1=2.175636829e-15 ub1=6.339562558e-19 lub1=-2.083859827e-24 pub1=7.703719778e-46 uc1=1.049519498e-10 luc1=-1.201922146e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.32 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.715915167e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.459526256e-9 k1=4.358592823e-01 lk1=7.071937821e-8 k2=-1.038961459e-03 lk2=-2.044280755e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.900741107e-01 ldsub=6.995323034e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.281156187e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.660463671e-9 nfactor=1.937174903e+00 lnfactor=4.667837382e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-1.179611964e-22 peta0=-2.602085214e-29 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.623763913e-02 lu0=-1.970509300e-9 ua=-1.360999372e-09 lua=-1.165401770e-16 ub=2.139076232e-18 lub=-6.698850589e-27 uc=7.394227196e-11 luc=9.320923477e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.773769876e+04 lvsat=5.786991954e-2 a0=4.059183813e-01 la0=5.474685953e-7 ags=1.104812894e+00 lags=3.982467176e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.707433317e-02 lketa=1.576549507e-8 dwg=0.0 dwb=0.0 pclm=1.378822570e+00 lpclm=-4.897940046e-7 pdiblc1=7.412342657e-01 lpdiblc1=-1.207114555e-7 pdiblc2=5.468089956e-03 lpdiblc2=-2.188954603e-9 pdiblcb=2.463605311e-02 lpdiblcb=-2.483743425e-08 wpdiblcb=-1.257674520e-23 ppdiblcb=7.589415207e-30 drout=-4.805786800e-01 ldrout=7.408682463e-07 pdrout=-2.220446049e-28 pscbe1=3.911445003e+07 lpscbe1=3.807402812e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.124887698e-06 lalpha0=3.184932520e-12 walpha0=6.352747104e-28 palpha0=1.588186776e-34 alpha1=1.292172822e+00 lalpha1=-2.212593006e-7 beta0=1.103727160e+01 lbeta0=3.493093664e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.306973693e-01 lkt1=-2.426211352e-8 kt2=-3.473922260e-02 lkt2=-1.092582431e-9 at=8.468137053e+04 lat=-1.905881962e-2 ute=-1.093884589e+00 lute=-7.964654023e-8 ua1=2.227271388e-09 lua1=-5.932625626e-16 ub1=-2.319771241e-18 lub1=8.710225781e-25 uc1=-8.247167459e-11 luc1=6.730469244e-17 puc1=2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.33 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.200522575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.978979228e-8 k1=3.751576387e-01 lk1=1.010939343e-7 k2=1.346271256e-02 lk2=-2.769931472e-08 pk2=-1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.588379951e-02 ldsub=1.220891243e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.337965066e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.817798513e-9 nfactor=2.559066539e+00 lnfactor=1.555947604e-7 eta0=0.49 etab=-0.000625 u0=2.996156444e-02 lu0=-3.833928011e-09 wu0=2.775557562e-23 ua=-1.106201234e-09 lua=-2.440388723e-16 ub=1.965615035e-18 lub=8.009957129e-26 uc=7.720017865e-11 luc=-6.981348409e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.193146463e+04 lvsat=2.074402684e-2 a0=1.5 ags=2.351090855e+00 lags=-5.838016037e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.120978342e-02 lketa=-2.180802844e-9 dwg=0.0 dwb=0.0 pclm=4.787930399e-01 lpclm=-3.942732802e-8 pdiblc1=8.451360799e-01 lpdiblc1=-1.727029882e-7 pdiblc2=-3.965600735e-04 lpdiblc2=7.456634899e-10 pdiblcb=1.753128000e-01 lpdiblcb=-1.002347223e-07 wpdiblcb=-5.551115123e-23 ppdiblcb=-4.163336342e-29 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.179906160e-06 lalpha0=3.007041669e-14 alpha1=0.85 beta0=1.690726552e+01 lbeta0=5.558015352e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.120971763e-01 lkt1=1.646961734e-8 kt2=-5.676512613e-02 lkt2=9.928981459e-09 wkt2=5.551115123e-23 at=7.053200633e+04 lat=-1.197860512e-02 wat=-5.820766091e-17 ute=-2.227083024e+00 lute=4.873957576e-7 ua1=-3.070875681e-10 lua1=6.749078496e-16 pua1=-4.135903063e-37 ub1=2.873772344e-19 lub1=-4.335710548e-25 pub1=1.925929944e-46 uc1=5.330152862e-11 luc1=-6.349964881e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.34 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.577424089e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.187966972e-09 wvth0=1.144804540e-07 pvth0=-2.866487536e-14 k1=4.486019531e-01 lk1=8.270413902e-8 k2=-1.722294551e-04 lk2=-2.428524795e-08 wk2=8.943928856e-08 pk2=-2.239479290e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.694175326e-01 ldsub=-7.410067063e-08 wdsub=7.083334704e-11 pdsub=-1.773603260e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.402784383e-02 lcdscd=-2.160334444e-9 cit=0.0 voff='-1.752724437e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.567402861e-09 wvoff=3.654943352e-07 pvoff=-9.151649209e-14 nfactor=3.427483312e+00 lnfactor=-6.184898374e-08 wnfactor=3.913900892e-06 pnfactor=-9.800055583e-13 eta0=1.750948185e+00 leta0=-3.157300771e-07 weta0=1.749325484e-14 peta0=-4.380153795e-21 etab=1.648869031e-01 letab=-4.144269092e-08 wetab=-1.027083532e-07 petab=2.571724727e-14 u0=-9.419103062e-03 lu0=6.026636707e-09 wu0=-2.927596720e-08 pu0=7.330438704e-15 ua=-4.113048799e-09 lua=5.088486964e-16 wua=-8.691280359e-16 pua=2.176218380e-22 ub=2.072514161e-18 lub=5.333299238e-26 wub=2.593446858e-24 pub=-6.493757522e-31 uc=2.240337191e-10 luc=-3.746393187e-17 wuc=-3.255036055e-16 puc=8.150317328e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.644436150e+05 lvsat=-2.245146301e-02 wvsat=-2.437154655e-01 pvsat=6.102415912e-8 a0=1.5 ags=-3.151405191e+00 lags=7.939738838e-07 wags=1.332267630e-21 pags=-1.249000903e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.285817898e-01 lketa=-9.226937466e-08 wketa=-9.916238423e-07 pketa=2.482936855e-13 dwg=0.0 dwb=0.0 pclm=-1.160773550e-02 lpclm=8.336461253e-08 wpclm=1.464414926e-06 ppclm=-3.666763177e-13 pdiblc1=-3.640440441e-01 lpdiblc1=1.300648323e-7 pdiblc2=-1.242883645e-02 lpdiblc2=3.758437203e-9 pdiblcb=-5.386335393e-01 lpdiblcb=7.853101555e-8 drout=2.279934293e+00 ldrout=-3.204840274e-7 pscbe1=8.221110918e+08 lpscbe1=-5.536418390e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.172683671e-05 lalpha0=-2.110004072e-12 alpha1=0.85 beta0=2.977423248e+01 lbeta0=-2.665971187e-06 wbeta0=5.592106345e-06 pbeta0=-1.400213100e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.851134190e-01 lkt1=-1.532597263e-08 wkt1=-1.433873422e-07 pkt1=3.590290000e-14 kt2=1.321436355e-02 lkt2=-7.593252940e-9 at=-1.878411818e+05 lat=5.271571582e-02 wat=2.150810133e-01 pat=-5.385434999e-8 ute=2.395681915e+00 lute=-6.701029782e-07 wute=8.881784197e-22 pute=-2.220446049e-28 ua1=8.604539016e-09 lua1=-1.556483242e-15 ub1=-6.989809769e-18 lub1=1.388571076e-24 uc1=-1.977121180e-10 luc1=6.221656150e-17 puc1=-2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.35 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='1.009711984e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-8.571921058e-08 wvth0=-9.526184081e-07 pvth0=1.638301555e-13 k1=0.90707349 k2=-6.968456304e-02 lk2=-1.174584859e-08 wk2=-1.591537790e-07 pk2=2.244915914e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587115367e-01 ldsub=-1.300531020e-11 wdsub=-1.652778098e-10 pdsub=2.485629509e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.333224414e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.418286027e-7 nfactor=-6.412814453e+00 lnfactor=1.713252170e-06 wnfactor=1.663312716e-05 pnfactor=-3.274439505e-12 eta0=6.941601366e-04 leta0=-3.211837743e-15 weta0=-4.081759674e-14 peta0=6.138599191e-21 etab=-6.485122645e-02 wetab=3.985556222e-8 u0=1.971647271e-02 lu0=7.708410583e-10 wu0=1.952747925e-08 pu0=-1.473263806e-15 ua=-1.243611304e-09 lua=-8.772002754e-18 wua=2.443222912e-16 pua=1.676542009e-23 ub=2.538334167e-18 lub=-3.069674433e-26 wub=-1.331608490e-24 pub=5.866890703e-32 uc=1.635189536e-11 wuc=1.263103613e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.428215842e+04 lvsat=3.323988799e-02 wvsat=4.467492978e-01 pvsat=-6.352946999e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.192202615e+00 lketa=1.820664449e-07 wketa=2.313788965e-06 pketa=-3.479730363e-13 dwg=0.0 dwb=0.0 pclm=1.847915313e+00 lpclm=-2.520766097e-07 wpclm=-3.239011085e-06 ppclm=4.817794038e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=2.068710412e+01 lbeta0=-1.026735016e-06 wbeta0=-1.304824814e-05 pbeta0=1.962339086e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.700731600e-01 wkt1=5.564087983e-8 kt2=-0.028878939 at=3.233014148e+05 lat=-3.948980831e-02 wat=-5.018556976e-01 pat=7.547458022e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.36 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.189614644e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.433377464e-8 k1=5.401372657e-01 lk1=2.266073161e-7 k2=-2.697132257e-02 lk2=-8.021815688e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.036636243e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.169372812e-8 nfactor=2.555062570e+00 lnfactor=-3.562583577e-7 eta0=0.08 etab=-0.07 u0=3.117200254e-02 lu0=-1.299030475e-8 ua=-7.258206658e-10 lua=4.388262947e-16 ub=1.538572798e-18 lub=-1.522285712e-24 uc=4.073563178e-11 luc=6.047391869e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.383068946e+00 la0=1.556811522e-6 ags=3.661934436e-01 lags=2.882567624e-7 a1=0.0 a2=0.42385546 b0=-5.268352994e-25 lb0=5.268373594e-29 b1=0.0 keta=-6.319216086e-03 lketa=1.322658029e-8 dwg=0.0 dwb=0.0 pclm=7.521971750e-02 lpclm=1.662288997e-7 pdiblc1=0.39 pdiblc2=3.376480374e-03 lpdiblc2=-1.827921882e-8 pdiblcb=5.966663033e-01 lpdiblcb=-6.216687341e-05 wpdiblcb=-3.330669074e-22 ppdiblcb=4.085620731e-26 drout=0.56 pscbe1=6.697834462e+08 lpscbe1=2.474695055e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.264150394e-01 lkt1=2.015047272e-07 wkt1=-4.440892099e-22 kt2=-4.662148499e-02 lkt2=1.111986337e-7 at=140000.0 ute=-1.907050456e+00 lute=2.335054779e-06 wute=3.552713679e-21 ua1=2.411546492e-10 lua1=1.794542099e-15 ub1=-5.160228553e-19 lub1=1.817292633e-24 wub1=7.703719778e-40 uc1=1.749183484e-11 luc1=-4.649096566e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.37 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.5216781+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.030982152 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.53725 eta0=0.08 etab=-0.07 u0=0.0305225 ua=-7.0387978e-10 ub=1.46246e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.460908 ags=0.380606 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.38 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.101977779e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.184706554e-8 k1=5.483118416e-01 lk1=2.524578124e-8 k2=-2.714422788e-02 lk2=-3.070489359e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077915297e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.634687659e-8 nfactor=2.613347438e+00 lnfactor=-6.088092565e-7 eta0=0.08 etab=-0.07 u0=3.032658085e-02 lu0=1.567429798e-9 ua=-7.552635323e-10 lua=4.110901092e-16 ub=1.520015626e-18 lub=-4.604675083e-25 uc=8.129900937e-11 luc=-8.262011279e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.583888020e+00 la0=-9.838882462e-7 ags=3.803559756e-01 lags=2.000293260e-9 a1=0.0 a2=0.42385546 b0=4.214805989e-24 lb0=-1.686087194e-29 b1=0.0 keta=-1.062994597e-02 lketa=3.977831183e-8 dwg=0.0 dwb=0.0 pclm=-3.218276199e-01 lpclm=3.243027455e-06 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=1.433768648e-03 lpdiblc2=8.230551467e-9 pdiblcb=-4.998476267e+00 lpdiblcb=1.989584970e-5 drout=0.56 pscbe1=7.870309262e+08 lpscbe1=5.188136624e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141197830e-01 lkt1=-1.776260414e-8 kt2=-3.996145347e-02 lkt2=-8.802098461e-9 at=140000.0 ute=-1.817602669e+00 lute=2.184320239e-7 ua1=3.751302750e-10 lua1=-3.540195022e-16 ub1=-4.995892647e-19 lub1=5.954632198e-25 uc1=3.182318579e-12 luc1=9.588479350e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.39 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.340087664e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.406198640e-9 k1=5.400936501e-01 lk1=5.812176032e-8 k2=-2.972741965e-02 lk2=-2.037111647e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064853034e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.112146062e-8 nfactor=2.121653639e+00 lnfactor=1.358158189e-6 eta0=0.08 etab=-0.07 u0=3.307966154e-02 lu0=-9.445969399e-9 ua=-5.124179691e-10 lua=-5.603870960e-16 ub=1.419962942e-18 lub=-6.021765480e-26 uc=5.718132279e-11 luc=1.386006354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.090729680e+00 la0=9.889379399e-7 ags=1.607499777e-01 lags=8.805101507e-7 a1=0.0 a2=0.42385546 b0=-2.107711977e-24 lb0=8.431672024e-30 b1=0.0 keta=-1.762043929e-03 lketa=4.303236316e-9 dwg=0.0 dwb=0.0 pclm=4.736370264e-01 lpclm=6.085784249e-8 pdiblc1=0.39 pdiblc2=2.133242770e-03 lpdiblc2=5.432381483e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.083402602e+08 lpscbe1=-3.336430185e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.149993040e-01 lkt1=-1.424417615e-8 kt2=-4.270927102e-02 lkt2=2.190246143e-9 at=1.649048680e+05 lat=-9.962920960e-2 ute=-1.940434682e+00 lute=7.098081038e-7 ua1=2.615718673e-11 lua1=1.042009300e-15 ub1=-2.936948702e-19 lub1=-2.281948629e-25 uc1=9.431295441e-12 luc1=7.088644271e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.40 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.885455964e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.753791758e-8 k1=6.317711558e-01 lk1=-1.252690968e-7 k2=-5.835540395e-02 lk2=3.689604566e-08 wk2=-1.110223025e-22 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.806460635e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.573495597e-8 nfactor=3.197578958e+00 lnfactor=-7.941131350e-7 eta0=1.574990403e-01 leta0=-1.550283827e-7 etab=-5.561937938e-02 letab=-2.876686407e-8 u0=3.244889907e-02 lu0=-8.184197843e-9 ua=-1.073516895e-10 lua=-1.370678036e-15 ub=6.470496747e-19 lub=1.485911089e-24 uc=5.334179128e-11 luc=2.154062782e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.441672627e+04 lvsat=-8.835179470e-3 a0=2.217278084e+00 la0=-1.264599349e-06 wa0=-3.552713679e-21 ags=5.700341213e-02 lags=1.088043847e-6 a1=0.0 a2=0.42385546 b0=4.215423954e-24 lb0=-4.217072185e-30 b1=0.0 keta=5.211352366e-02 lketa=-1.034689642e-07 wketa=2.602085214e-23 pketa=1.474514955e-29 dwg=0.0 dwb=0.0 pclm=1.187494024e-01 lpclm=7.707718516e-7 pdiblc1=1.593398571e-01 lpdiblc1=4.614104738e-7 pdiblc2=6.418427744e-03 lpdiblc2=-3.139663973e-9 pdiblcb=-4.981802656e-02 lpdiblcb=4.964575696e-8 drout=8.601173000e-01 ldrout=-6.003519459e-7 pscbe1=1.163762255e+09 lpscbe1=-7.443472606e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.188739200e-09 lalpha0=5.763378680e-14 alpha1=6.289135890e-01 lalpha1=4.422592668e-7 beta0=1.319073842e+01 lbeta0=1.338784839e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.893162635e-01 lkt1=1.344188007e-7 kt2=-4.739960715e-02 lkt2=1.157275232e-8 at=1.645893428e+05 lat=-9.899803587e-2 ute=-1.997861131e+00 lute=8.246834563e-7 ua1=-5.405457877e-10 lua1=2.175636829e-15 ub1=6.339562558e-19 lub1=-2.083859827e-24 pub1=1.540743956e-45 uc1=1.049519498e-10 luc1=-1.201922146e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.41 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.715915167e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.459526256e-9 k1=4.358592823e-01 lk1=7.071937821e-8 k2=-1.038961459e-03 lk2=-2.044280755e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.900741107e-01 ldsub=6.995323034e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.281156187e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.660463671e-9 nfactor=1.937174903e+00 lnfactor=4.667837382e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=6.938893904e-23 peta0=-3.018418848e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.623763913e-02 lu0=-1.970509300e-9 ua=-1.360999372e-09 lua=-1.165401770e-16 ub=2.139076232e-18 lub=-6.698850589e-27 uc=7.394227196e-11 luc=9.320923477e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.773769876e+04 lvsat=5.786991954e-2 a0=4.059183813e-01 la0=5.474685953e-7 ags=1.104812894e+00 lags=3.982467176e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.707433317e-02 lketa=1.576549507e-8 dwg=0.0 dwb=0.0 pclm=1.378822570e+00 lpclm=-4.897940046e-7 pdiblc1=7.412342657e-01 lpdiblc1=-1.207114555e-7 pdiblc2=5.468089956e-03 lpdiblc2=-2.188954603e-09 ppdiblc2=3.469446952e-30 pdiblcb=2.463605311e-02 lpdiblcb=-2.483743425e-08 wpdiblcb=-5.204170428e-24 ppdiblcb=-3.686287386e-30 drout=-4.805786800e-01 ldrout=7.408682463e-07 pdrout=-4.440892099e-28 pscbe1=3.911445003e+07 lpscbe1=3.807402812e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.124887698e-06 lalpha0=3.184932520e-12 walpha0=-2.117582368e-28 palpha0=-1.588186776e-33 alpha1=1.292172822e+00 lalpha1=-2.212593006e-7 beta0=1.103727160e+01 lbeta0=3.493093664e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.306973693e-01 lkt1=-2.426211352e-8 kt2=-3.473922260e-02 lkt2=-1.092582431e-9 at=8.468137053e+04 lat=-1.905881962e-2 ute=-1.093884589e+00 lute=-7.964654023e-8 ua1=2.227271388e-09 lua1=-5.932625626e-16 ub1=-2.319771241e-18 lub1=8.710225781e-25 pub1=1.540743956e-45 uc1=-8.247167459e-11 luc1=6.730469244e-17 puc1=2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.42 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.200522575e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.978979228e-8 k1=3.751576387e-01 lk1=1.010939343e-7 k2=1.346271256e-02 lk2=-2.769931472e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.588379951e-02 ldsub=1.220891243e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.337965066e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.817798513e-9 nfactor=2.559066539e+00 lnfactor=1.555947604e-7 eta0=0.49 etab=-0.000625 u0=2.996156444e-02 lu0=-3.833928011e-9 ua=-1.106201234e-09 lua=-2.440388723e-16 ub=1.965615035e-18 lub=8.009957129e-26 uc=7.720017865e-11 luc=-6.981348409e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.193146463e+04 lvsat=2.074402684e-2 a0=1.5 ags=2.351090855e+00 lags=-5.838016037e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.120978342e-02 lketa=-2.180802844e-9 dwg=0.0 dwb=0.0 pclm=4.787930399e-01 lpclm=-3.942732802e-8 pdiblc1=8.451360799e-01 lpdiblc1=-1.727029882e-7 pdiblc2=-3.965600735e-04 lpdiblc2=7.456634899e-10 pdiblcb=1.753128000e-01 lpdiblcb=-1.002347223e-07 ppdiblcb=-2.775557562e-29 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.179906160e-06 lalpha0=3.007041669e-14 alpha1=0.85 beta0=1.690726552e+01 lbeta0=5.558015352e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.120971763e-01 lkt1=1.646961734e-8 kt2=-5.676512613e-02 lkt2=9.928981459e-9 at=7.053200633e+04 lat=-1.197860512e-02 wat=-1.164153218e-16 ute=-2.227083024e+00 lute=4.873957576e-07 wute=3.552713679e-21 ua1=-3.070875681e-10 lua1=6.749078496e-16 ub1=2.873772344e-19 lub1=-4.335710548e-25 pub1=3.851859889e-46 uc1=5.330152862e-11 luc1=-6.349964881e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.43 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='7.130707622e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.308078869e-08 wvth0=-1.823896187e-07 pvth0=4.566871902e-14 k1=4.486019531e-01 lk1=8.270413902e-8 k2=1.044049621e-01 lk2=-5.047043552e-08 wk2=-1.104330322e-07 pk2=2.765143736e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.694545940e-01 ldsub=-7.410995047e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.402784383e-02 lcdscd=-2.160334444e-9 cit=0.0 voff='1.596149487e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.031585425e-8 nfactor=-4.621753268e-01 lnfactor=9.120865325e-07 wnfactor=1.134797985e-05 pnfactor=-2.841432022e-12 eta0=1.750948194e+00 leta0=-3.157300794e-7 etab=1.111478406e-01 letab=-2.798691333e-08 wetab=-5.204170428e-23 petab=-9.540979118e-30 u0=-4.060307077e-02 lu0=1.383482156e-08 wu0=3.032414160e-08 pu0=-7.592892140e-15 ua=-4.200311338e-09 lua=5.306984508e-16 wua=-7.023482067e-16 pua=1.758616698e-22 ub=1.810468165e-18 lub=1.189469512e-25 wub=3.094280170e-24 pub=-7.747799061e-31 uc=-1.786936147e-10 luc=6.337536798e-17 wuc=4.442057895e-16 puc=-1.112251318e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.705393572e+05 lvsat=1.061318002e-03 wvsat=-6.424170402e-02 pvsat=1.608554451e-8 a0=1.5 ags=-3.151405191e+00 lags=7.939738838e-07 wags=1.110223025e-21 pags=-4.440892099e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.262738469e-01 lketa=9.673968308e-08 wketa=4.510879545e-07 pketa=-1.129483640e-13 dwg=0.0 dwb=0.0 pclm=5.974971298e-01 lpclm=-6.914976379e-08 wpclm=3.002681248e-07 ppclm=-7.518443603e-14 pdiblc1=-3.640440441e-01 lpdiblc1=1.300648323e-07 ppdiblc1=1.110223025e-28 pdiblc2=-1.242883645e-02 lpdiblc2=3.758437203e-09 ppdiblc2=-3.469446952e-30 pdiblcb=-5.386335393e-01 lpdiblcb=7.853101555e-8 drout=2.279934293e+00 ldrout=-3.204840274e-7 pscbe1=8.221110918e+08 lpscbe1=-5.536418390e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.172683671e-05 lalpha0=-2.110004072e-12 alpha1=0.85 beta0=3.218755257e+01 lbeta0=-3.270244819e-06 wbeta0=9.796676176e-07 pbeta0=-2.452999544e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.845705887e-03 lkt1=-6.071377660e-08 wkt1=-4.898338088e-07 pkt1=1.226499772e-13 kt2=1.321436355e-02 lkt2=-7.593252940e-9 at=-7.530649842e+04 lat=2.453804393e-2 ute=2.395681915e+00 lute=-6.701029782e-07 wute=-1.776356839e-21 pute=2.220446049e-28 ua1=8.604539016e-09 lua1=-1.556483242e-15 ub1=-6.989809769e-18 lub1=1.388571076e-24 wub1=6.162975822e-39 uc1=-1.977121180e-10 luc1=6.221656150e-17 wuc1=-2.067951531e-31 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.44 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.742518151e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=7.077555593e-8 k1=0.90707349 k2=-1.753785943e-01 wk2=4.285309275e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=4.593988963e+00 wnfactor=-4.403537812e-6 eta0=0.00069413878 etab=-0.043998 u0=3.609045366e-02 wu0=-1.176716085e-8 ua=-1.258377146e-09 wua=2.725433889e-16 ub=2.469852232e-18 wub=-1.200722940e-24 uc=1.726286130e-10 wuc=-1.723722651e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.764227882e+05 wvsat=2.492873415e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.100039224e-01 wketa=-1.750428614e-7 dwg=0.0 dwb=0.0 pclm=2.141644591e-01 wpclm=-1.165178348e-7 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.405890525e+01 wbeta0=-3.801560678e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.404133650e-01 wkt1=1.900780339e-7 kt2=-0.028878939 at=60720.487 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.45 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.147606461e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.316470859e-07 wvth0=6.684518484e-09 pvth0=2.959405566e-13 k1=4.541949221e-01 lk1=6.293191300e-06 wk1=1.367550666e-07 pk1=-9.653403231e-12 k2=7.007422791e-03 lk2=-2.583315143e-06 wk2=-5.406840672e-08 pk2=3.983033054e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.018026242e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.372768656e-07 wvoff=-2.961301678e-09 pvoff=-4.439097255e-13 nfactor=3.031445903e+00 lnfactor=-4.402090560e-05 wnfactor=-7.580411676e-07 pnfactor=6.948102061e-11 eta0=0.08 etab=-0.07 u0=3.067418663e-02 lu0=1.816914148e-07 wu0=7.921455833e-10 pu0=-3.097857288e-13 ua=-7.553503436e-10 lua=-1.503068083e-15 wua=4.698886358e-17 pua=3.090023894e-21 ub=1.573902636e-18 lub=1.192500338e-23 wub=-5.621832226e-26 pub=-2.139789120e-29 uc=-7.507744370e-11 luc=5.440548323e-15 wuc=1.842866298e-16 puc=-7.694942602e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.115597269e+00 la0=1.093868004e-05 wa0=4.256121660e-07 pa0=-1.492882322e-11 ags=2.935003530e-01 lags=4.342243523e-06 wags=1.156722990e-07 pags=-6.450874000e-12 a1=0.0 a2=0.42385546 b0=-9.341743695e-24 lb0=3.465189942e-28 wb0=1.402665247e-29 pb0=-4.675630041e-34 b1=0.0 keta=-5.287854826e-03 lketa=-2.374454108e-07 wketa=-1.641145353e-09 pketa=3.988798004e-13 dwg=0.0 dwb=0.0 pclm=5.204228147e-02 lpclm=6.297866827e-07 wpclm=3.688090967e-08 ppclm=-7.376326138e-13 pdiblc1=0.39 pdiblc2=6.404713417e-03 lpdiblc2=-1.172087523e-07 wpdiblc2=-4.818651604e-09 ppdiblc2=1.574208287e-13 pdiblcb=9.468965799e+00 lpdiblcb=-2.559619141e-04 wpdiblcb=-1.411797559e-05 ppdiblcb=3.083748081e-10 drout=0.56 pscbe1=3.024234342e+08 lpscbe1=1.160693397e+04 wpscbe1=5.845586803e+02 ppscbe1=-1.453160212e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.378762636e-01 lkt1=-9.000463289e-07 wkt1=1.823758136e-08 pkt1=1.752834306e-12 kt2=-4.788606706e-02 lkt2=-1.002704226e-06 wkt2=2.012256105e-09 pkt2=1.772489014e-12 at=140000.0 ute=-1.882225704e+00 lute=-2.619372321e-05 wute=-3.950218955e-08 pute=4.539618974e-11 ua1=7.039615771e-10 lua1=-6.450349343e-14 wua1=-7.364378216e-16 pua1=1.054962186e-19 ub1=-1.129782614e-18 lub1=4.292257663e-23 wub1=9.766403063e-25 pub1=-6.540845432e-29 uc1=-3.617304502e-12 luc1=2.583013194e-15 wuc1=3.358974910e-17 puc1=-4.184177458e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.46 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.081784205e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.148125704e-8 k1=7.688483357e-01 wk1=-3.459056589e-7 k2=-1.221558092e-01 wk2=1.450793527e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.993901280e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-2.515635404e-8 nfactor=8.304436521e-01 wnfactor=2.715941947e-6 eta0=0.08 etab=-0.07 u0=3.975857977e-02 wu0=-1.469683805e-8 ua=-8.305022785e-10 wua=2.014870378e-16 ub=2.170141148e-18 wub=-1.126091966e-24 uc=1.969446544e-10 wuc=-2.004529786e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.662520578e+00 wa0=-3.208144023e-7 ags=5.106082847e-01 wags=-2.068650954e-7 a1=0.0 a2=0.42385546 b0=7.983867301e-24 wb0=-9.351040706e-30 b1=0.0 keta=-1.715989327e-02 wketa=1.830245477e-8 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=5.443903725e-04 wpdiblc2=3.052235953e-9 pdiblcb=-3.328879708e+00 wpdiblcb=1.300463382e-6 drout=0.56 pscbe1=8.827587873e+08 wpscbe1=-1.420072214e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.828777003e-01 wkt1=1.058775833e-7 kt2=-9.802029824e-02 wkt2=9.063497424e-8 at=140000.0 ute=-3.191886260e+00 wute=2.230262924e-6 ua1=-2.521150043e-09 wua1=4.538269990e-15 ub1=1.016304261e-18 wub1=-2.293718474e-24 uc1=1.255308304e-10 wuc1=-1.756150339e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.47 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.883647337e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.585172418e-07 wvth0=3.474165700e-08 pvth0=-1.060883846e-13 k1=8.035721491e-01 lk1=-2.778040849e-07 wk1=-4.061809223e-07 pk1=4.822256752e-13 k2=-1.328439994e-01 lk2=8.550970015e-08 wk2=1.681939158e-07 pk2=-1.849255426e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.259995804e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.871530767e-08 wvoff=-4.008588688e-08 pvoff=1.194421002e-13 nfactor=5.403248505e-01 lnfactor=2.321063849e-06 wnfactor=3.298680608e-06 pnfactor=-4.662137141e-12 eta0=0.08 etab=-0.07 u0=3.760175408e-02 lu0=1.725544884e-08 wu0=-1.157656120e-08 pu0=-2.496343480e-14 ua=-1.131328124e-09 lua=2.406724389e-15 wua=5.984097735e-16 pua=-3.175537082e-21 ub=2.406384417e-18 lub=-1.890038523e-24 wub=-1.410427249e-24 pub=2.274793440e-30 uc=2.348933654e-10 luc=-3.036045256e-16 wuc=-2.444057903e-16 puc=3.516396790e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.795072254e+00 la0=-1.060465236e-06 wa0=-3.360452231e-07 pa0=1.218525220e-13 ags=4.741605558e-01 lags=2.915960822e-07 wags=-1.492657878e-07 pags=-4.608169823e-13 a1=0.0 a2=0.42385546 b0=1.596851503e-23 lb0=-6.388030379e-29 wb0=-1.870299548e-29 pb0=7.481929478e-35 b1=0.0 keta=-4.500597978e-03 lketa=-1.012793121e-07 wketa=-9.753275958e-09 pketa=2.244568156e-13 dwg=0.0 dwb=0.0 pclm=-1.982495104e-01 lpclm=2.254354259e-06 wpclm=-1.966426782e-07 ppclm=1.573218313e-12 pdiblc1=0.39 pdiblc2=-2.811470661e-03 lpdiblc2=2.684820041e-08 wpdiblc2=6.755203088e-09 ppdiblc2=-2.962518494e-14 pdiblcb=-6.633082370e+00 lpdiblcb=2.643491324e-05 wpdiblcb=2.601053884e-06 ppdiblcb=-1.040523255e-11 drout=0.56 pscbe1=8.127710168e+08 lpscbe1=5.599295292e+02 wpscbe1=-4.095871327e+01 ppscbe1=-8.084275750e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.778964287e-01 lkt1=-3.985212037e-08 wkt1=1.014840773e-07 pkt1=3.514976597e-14 kt2=-9.402411438e-02 lkt2=-3.197103339e-08 wkt2=8.602677667e-08 pkt2=3.686738236e-14 at=140000.0 ute=-2.731402619e+00 lute=-3.684049175e-06 wute=1.454076861e-06 pute=6.209791988e-12 ua1=-2.069306895e-09 lua1=-3.614921859e-15 wua1=3.889691091e-15 pua1=5.188884788e-21 ub1=7.169968903e-19 lub1=2.394575999e-24 wub1=-1.935882986e-24 pub1=-2.862823816e-30 uc1=9.720168463e-11 luc1=2.266442426e-16 wuc1=-1.496075641e-16 puc1=-2.080699273e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.48 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.027525303e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.990786706e-07 wvth0=-1.093879644e-07 pvth0=4.704864557e-13 k1=8.162252253e-01 lk1=-3.284213370e-07 wk1=-4.393921600e-07 pk1=6.150836112e-13 k2=-1.634676523e-01 lk2=2.080162859e-07 wk2=2.128130753e-07 pk2=-3.634196270e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.631427178e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.634872234e-07 wvoff=9.015565734e-08 pvoff=-4.015750011e-13 nfactor=-1.788857713e+00 lnfactor=1.163870481e-05 wnfactor=6.222569905e-06 pnfactor=-1.635883757e-11 eta0=0.08 etab=-0.07 u0=4.552714092e-02 lu0=-1.444919734e-08 wu0=-1.980695199e-08 pu0=7.961346428e-15 ua=-1.267105727e-09 lua=2.949887889e-15 wua=1.200890858e-15 pua=-5.585696988e-21 ub=3.455159251e-18 lub=-6.085547930e-24 wub=-3.238489845e-24 pub=9.587758597e-30 uc=2.259710626e-10 luc=-2.679118256e-16 wuc=-2.685853231e-16 puc=4.483672644e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=-7.819323836e-02 la0=6.433329182e-06 wa0=1.860039242e-06 pa0=-8.663344008e-12 ags=2.261714747e-01 lags=1.283649370e-06 wags=-1.041014338e-07 pags=-6.414920578e-13 a1=0.0 a2=0.42385546 b0=-7.985428147e-24 lb0=3.194483489e-29 wb0=9.352868834e-30 pb0=-3.741513231e-35 b1=0.0 keta=-8.578170914e-02 lketa=2.238769134e-07 wketa=1.336956201e-07 pketa=-3.493948571e-13 dwg=0.0 dwb=0.0 pclm=3.743929643e-01 lpclm=-3.643954289e-08 wpclm=1.579213199e-07 ppclm=1.548236861e-13 pdiblc1=0.39 pdiblc2=4.200365935e-03 lpdiblc2=-1.201887603e-09 wpdiblc2=-3.289293199e-09 ppdiblc2=1.055672761e-14 pdiblcb=-0.025 drout=0.56 pscbe1=1.137107800e+09 lpscbe1=-7.375444211e+02 wpscbe1=-5.231487183e+02 ppscbe1=1.120520981e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.687060681e-01 lkt1=-7.661715600e-08 wkt1=8.546045877e-08 pkt1=9.925050520e-14 kt2=-9.572389649e-02 lkt2=-2.517124032e-08 wkt2=8.435909867e-08 pkt2=4.353874644e-14 at=1.540269232e+05 lat=-5.611317715e-02 wat=1.730944263e-02 pat=-6.924453851e-8 ute=-2.475232310e+00 lute=-4.708830573e-06 wute=8.509924483e-07 pute=8.622365445e-12 ua1=2.051509368e-09 lua1=-2.009979815e-14 wua1=-3.222825455e-15 pua1=3.364173197e-20 ub1=-3.455223968e-18 lub1=1.908509077e-23 wub1=5.030757885e-24 pub1=-3.073211126e-29 uc1=5.343414689e-11 luc1=4.017315067e-16 wuc1=-7.001918534e-17 puc1=-5.264545613e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.49 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='3.687347598e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.690483714e-07 wvth0=1.906480352e-07 pvth0=-1.297028576e-13 k1=7.214844871e-01 lk1=-1.389028168e-07 wk1=-1.427556207e-07 pk1=2.169454788e-14 k2=-7.886381423e-02 lk2=3.877552962e-08 wk2=3.263384380e-08 pk2=-2.990713817e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.195885626e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.067882993e-07 wvoff=-1.432491147e-07 pvoff=6.532580418e-14 nfactor=4.291614130e+00 lnfactor=-5.246163369e-07 wnfactor=-1.740874715e-06 pnfactor=-4.288346240e-13 eta0=1.574991798e-01 leta0=-1.550286617e-07 weta0=-2.219593073e-13 peta0=4.440054006e-19 etab=-5.561937938e-02 letab=-2.876686407e-8 u0=4.683292755e-02 lu0=-1.706128116e-08 wu0=-2.288847024e-08 pu0=1.412558781e-14 ua=2.155401034e-09 lua=-3.896463832e-15 wua=-3.600587169e-15 pua=4.019136442e-21 ub=-1.869282507e-18 lub=4.565417444e-24 wub=4.004093454e-24 pub=-4.900239851e-30 uc=9.601980517e-11 luc=-7.958499875e-18 wuc=-6.791104819e-17 puc=4.694025095e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.246311426e+05 lvsat=-8.927973597e-02 wvsat=-6.399086828e-02 pvsat=1.280067570e-7 a0=4.526685794e+00 la0=-2.778229392e-06 wa0=-3.674826544e-06 pa0=2.408551696e-12 ags=-7.321951340e-01 lags=3.200757309e-06 wags=1.255805873e-06 pags=-3.361838395e-12 a1=0.0 a2=0.42385546 b0=1.597085629e-23 lb0=-1.597710090e-29 wb0=-1.870573767e-29 pb0=1.871305161e-35 b1=0.0 keta=2.733848571e-01 lketa=-4.945966531e-07 wketa=-3.520962391e-07 pketa=6.223788059e-13 dwg=0.0 dwb=0.0 pclm=-7.375659547e-01 lpclm=2.187913071e-06 wpclm=1.362604961e-06 ppclm=-2.255014628e-12 pdiblc1=-6.269973846e-01 lpdiblc1=2.034392415e-06 wpdiblc1=1.251252845e-06 ppdiblc1=-2.502994930e-12 pdiblc2=1.096807117e-02 lpdiblc2=-1.473994425e-08 wpdiblc2=-7.239583709e-09 ppdiblc2=1.845885319e-14 pdiblcb=-1.870209292e-01 lpdiblcb=3.241052085e-07 wpdiblcb=2.183230212e-07 ppdiblcb=-4.367314066e-13 drout=1.243151065e+00 ldrout=-1.366569242e-06 wdrout=-6.094994142e-07 pdrout=1.219237143e-12 pscbe1=2.178175661e+09 lpscbe1=-2.820087199e+03 wpscbe1=-1.614177217e+03 ppscbe1=3.303004571e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.250411477e-08 lalpha0=2.250522187e-13 walpha0=1.331755843e-13 palpha0=-2.664032403e-19 alpha1=-4.144573239e-01 lalpha1=2.529409051e-06 walpha1=1.660255618e-06 palpha1=-3.321160396e-12 beta0=1.132438778e+01 lbeta0=5.072215870e-06 wbeta0=2.969815531e-06 pbeta0=-5.940792260e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-5.638384684e-01 lkt1=3.137239412e-07 wkt1=2.777070624e-07 pkt1=-2.853178704e-13 kt2=-1.819142678e-01 lkt2=1.472432028e-07 wkt2=2.140453777e-07 pkt2=-2.158845190e-13 at=2.423775981e+05 lat=-2.328490721e-01 wat=-1.237799390e-01 pat=2.129893906e-7 ute=-8.132841351e+00 lute=6.608599634e-06 wute=9.762238195e-06 pute=-9.203610346e-12 ua1=-1.871311911e-08 lua1=2.143757777e-14 wua1=2.891696191e-14 pua1=-3.065040943e-20 ub1=1.552380502e-17 lub1=-1.888038801e-23 wub1=-2.369335273e-23 pub1=2.672734110e-29 uc1=6.165518829e-10 luc1=-7.247241445e-16 wuc1=-8.140793008e-16 puc1=9.619565972e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.50 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.139550910e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.377125911e-08 wvth0=9.171350142e-08 pvth0=-3.072964041e-14 k1=5.498563303e-01 lk1=3.279244655e-08 wk1=-1.813968907e-07 pk1=6.035092660e-14 k2=-2.237087615e-02 lk2=-1.773949720e-08 wk2=3.394423860e-08 pk2=-4.301620980e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.439825452e-01 ldsub=1.160628176e-07 wdsub=7.334283483e-08 pdsub=-7.337151188e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.688400371e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.791852179e-08 wvoff=-1.292591575e-07 pvoff=5.133037692e-14 nfactor=5.262818723e+00 lnfactor=-1.496200671e-06 wnfactor=-5.291904123e-06 pnfactor=3.123583237e-12 eta0=-4.853189795e-01 leta0=4.880408395e-07 weta0=4.439186145e-13 peta0=-2.221328794e-19 etab=-1.673183512e-01 letab=8.297578205e-08 wetab=-1.387787871e-09 petab=1.388330496e-15 u0=3.342368152e-02 lu0=-3.646792113e-09 wu0=-1.143473246e-08 pu0=2.667371616e-15 ua=-1.572391840e-09 lua=-1.672133912e-16 wua=3.363765737e-16 pua=8.063334670e-23 ub=2.416742957e-18 lub=2.777161436e-25 wub=-4.418349549e-25 pub=-4.525730843e-31 uc=1.051755471e-10 luc=-1.711782169e-17 wuc=-4.969969919e-17 puc=2.872178131e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.222711279e+04 lvsat=8.764767099e-02 wvsat=1.113309466e-01 pvsat=-4.738360877e-8 a0=1.999279674e+00 la0=-2.498350552e-07 wa0=-2.535423410e-06 pa0=1.268703055e-12 ags=3.502281559e+00 lags=-1.035375064e-06 wags=-3.814952834e-06 pags=1.710902979e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.956634428e-01 lketa=1.747132447e-07 wketa=5.228647920e-07 pketa=-2.529243350e-13 dwg=0.0 dwb=0.0 pclm=2.778889873e+00 lpclm=-1.329917691e-06 wpclm=-2.227845895e-06 ppclm=1.336840095e-12 pdiblc1=1.315115923e+00 lpdiblc1=9.151974087e-08 wpdiblc1=-9.131845967e-07 ppdiblc1=-3.377111933e-13 pdiblc2=-7.200110974e-03 lpdiblc2=3.435341654e-09 wpdiblc2=2.015817339e-08 ppdiblc2=-8.949616425e-15 pdiblcb=2.990418583e-01 lpdiblcb=-1.621476295e-07 wpdiblcb=-4.366460423e-07 ppdiblcb=2.184937498e-13 drout=-1.246646210e+00 ldrout=1.124201544e-06 wdrout=1.218998828e-06 pdrout=-6.099760428e-13 pscbe1=-2.082745344e+09 lpscbe1=1.442499825e+03 wpscbe1=3.376392422e+03 ppscbe1=-1.689516380e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.191613745e-05 lalpha0=1.206331251e-11 walpha0=1.398900585e-11 palpha0=-1.412765113e-17 alpha1=3.378914648e+00 lalpha1=-1.265446129e-06 walpha1=-3.320511236e-06 palpha1=1.661553938e-12 beta0=3.165609568e+00 lbeta0=1.323418416e-05 wbeta0=1.252571924e-05 pbeta0=-1.550043233e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.977656780e-01 lkt1=-5.249198363e-08 wkt1=-5.240229027e-08 pkt1=4.492055498e-14 kt2=-3.093520178e-02 lkt2=-3.794896065e-09 wkt2=-6.053117709e-09 pkt2=4.300034952e-15 at=-1.751247404e+04 lat=2.714261702e-02 wat=1.626151376e-01 pat=-7.351766643e-8 ute=-1.725156088e+00 lute=1.984089653e-07 wute=1.004505722e-06 pute=-4.424535988e-13 ua1=4.536754493e-09 lua1=-1.821386531e-15 wua1=-3.674946516e-15 pua1=1.954242440e-21 ub1=-6.402392183e-18 lub1=3.054382338e-24 wub1=6.496437912e-24 pub1=-3.474253751e-30 uc1=-3.037441950e-10 luc1=1.959317693e-16 wuc1=3.520981280e-16 puc1=-2.046768070e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.51 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.108066580e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.469239337e-08 wvth0=1.471198627e-08 pvth0=7.801224758e-15 k1=8.096097127e-01 lk1=-9.718580823e-08 wk1=-6.913183872e-07 pk1=3.155110541e-13 k2=-1.525537672e-01 lk2=4.740284985e-08 wk2=2.641723953e-07 pk2=-1.195057185e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.427064753e-01 ldsub=2.595194233e-07 wdsub=3.637424462e-07 pdsub=-2.186848638e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-3.951074185e-03 lcdscd=4.679193362e-09 wcdscd=1.487982199e-08 pcdscd=-7.445729005e-15 cit=0.0 voff='-1.936092737e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.550148279e-08 wvoff=9.517658724e-08 pvoff=-6.097524982e-14 nfactor=-2.102127371e+00 lnfactor=2.189152070e-06 wnfactor=7.417087520e-06 pnfactor=-3.235881801e-12 eta0=-8.766473704e-01 leta0=6.838580443e-07 weta0=2.174666695e-06 peta0=-1.088183642e-12 etab=-1.235114990e-01 letab=6.105522749e-08 wetab=1.955421585e-07 petab=-9.715364230e-14 u0=4.938501893e-02 lu0=-1.163370170e-08 wu0=-3.090741656e-08 pu0=1.241132749e-14 ua=9.766524450e-10 lua=-1.442732210e-15 wua=-3.314324254e-15 pua=1.907411184e-21 ub=5.501094211e-19 lub=1.211762766e-24 wub=2.252411985e-24 pub=-1.800750005e-30 uc=1.182038829e-10 luc=-2.363708366e-17 wuc=-6.524681633e-17 puc=3.650141880e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.782240369e+04 lvsat=1.256424339e-02 wvsat=-9.373909655e-03 pvsat=1.301601498e-8 a0=1.5 ags=6.285719295e+00 lags=-2.428182256e-06 wags=-6.260946028e-06 pags=2.934855959e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.738498956e-01 lketa=6.371974195e-08 wketa=2.269749373e-07 pketa=-1.048637147e-13 dwg=0.0 dwb=0.0 pclm=-3.105287977e-01 lpclm=2.159996071e-07 wpclm=1.256002060e-06 ppclm=-4.064460672e-13 pdiblc1=3.405711364e+00 lpdiblc1=-9.545954024e-07 wpdiblc1=-4.074494937e-06 ppdiblc1=1.244180049e-12 pdiblc2=1.301292123e-02 lpdiblc2=-6.679077745e-09 wpdiblc2=-2.133772985e-08 ppdiblc2=1.181456009e-14 pdiblcb=5.152367198e-01 lpdiblcb=-2.703295924e-07 wpdiblcb=-5.409012179e-07 ppdiblcb=2.706621013e-13 drout=-3.872249845e-01 ldrout=6.941548972e-07 wdrout=2.207410659e-06 pdrout=-1.104568427e-12 pscbe1=7.760354425e+08 lpscbe1=1.199164891e+01 wpscbe1=3.813341047e+01 ppscbe1=-1.908161540e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.194049799e-05 lalpha0=1.256668402e-13 walpha0=-1.394022167e-11 palpha0=-1.521170442e-19 alpha1=0.85 beta0=2.668988296e+01 lbeta0=1.462849472e-06 wbeta0=-1.556651174e-05 pbeta0=-1.443332773e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.441287665e-01 lkt1=2.074678861e-08 wkt1=5.097001168e-08 pkt1=-6.806014564e-15 kt2=-9.282801876e-02 lkt2=2.717571252e-08 wkt2=5.738478941e-08 pkt2=-2.744372283e-14 at=6.762685837e+04 lat=-1.546033867e-02 wat=4.622793453e-03 pat=5.540280664e-9 ute=-5.278952689e+00 lute=1.976696800e-06 wute=4.856263190e-06 pute=-2.369838370e-12 ua1=-7.334290857e-09 lua1=4.118777723e-15 wua1=1.118198102e-14 pua1=-5.480030385e-21 ub1=6.859661847e-18 lub1=-3.581830140e-24 wub1=-1.045809531e-23 pub1=5.009642083e-30 uc1=3.942250277e-10 luc1=-1.533257481e-16 wuc1=-5.424917905e-16 puc1=2.429679369e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.52 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.376189068e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.366839159e-09 wvth0=9.679674262e-08 pvth0=-1.275205947e-14 k1=-8.299245227e-01 lk1=3.133388085e-07 wk1=2.034445026e-06 pk1=-3.669955728e-13 k2=5.216452548e-01 lk2=-1.214105175e-07 wk2=-7.743633100e-07 pk2=1.405342752e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.015073901e+00 ldsub=-2.807693628e-07 wdsub=-1.822957556e-06 pdsub=3.288451366e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=4.742453735e-02 lcdscd=-8.184797384e-09 wcdscd=-5.314222139e-08 pcdscd=9.586378458e-15 cit=0.0 voff='3.494286767e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.004703326e-07 wvoff=-5.306269853e-07 pvoff=9.572033250e-14 nfactor=2.037870997e+01 lnfactor=-3.439847272e-06 wnfactor=-2.181491215e-05 pnfactor=4.083547828e-12 eta0=6.631831660e+00 leta0=-1.196197529e-06 weta0=-7.766666768e-06 peta0=1.401036785e-12 etab=5.437986136e-01 letab=-1.060332189e-07 wetab=-6.884520813e-07 petab=1.241905594e-13 u0=-7.188802152e-02 lu0=1.873197617e-08 wu0=8.010606922e-08 pu0=-1.538545023e-14 ua=-1.481374604e-08 lua=2.511041456e-15 wua=1.618619485e-14 pua=-2.975343294e-21 ub=1.711800486e-17 lub=-2.936689142e-24 wub=-2.126371514e-23 pub=4.087476583e-30 uc=3.958479684e-11 luc=-3.951572089e-18 wuc=9.687201329e-17 puc=-4.091677066e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.665296006e+05 lvsat=-4.639420366e-03 wvsat=-5.786121094e-02 pvsat=2.515679883e-8 a0=1.5 ags=-1.542547809e+01 lags=3.008106169e-06 wags=1.953102031e-05 pags=-3.523220285e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.884184678e-01 lketa=-5.202809583e-08 wketa=-6.861604738e-07 pketa=1.237771740e-13 dwg=0.0 dwb=0.0 pclm=1.611738334e+00 lpclm=-2.653187824e-07 wpclm=-1.313635078e-06 ppclm=2.369679454e-13 pdiblc1=-2.374721304e+00 lpdiblc1=4.927729139e-07 wpdiblc1=3.199474105e-06 ppdiblc1=-5.771563332e-13 pdiblc2=-7.053066217e-02 lpdiblc2=1.423948365e-08 wpdiblc2=9.245406537e-08 ppdiblc2=-1.667788131e-14 pdiblcb=-1.752647538e+00 lpdiblcb=2.975282149e-07 wpdiblcb=1.931790064e-06 ppdiblcb=-3.484775414e-13 drout=7.234309237e+00 ldrout=-1.214208678e-06 wdrout=-7.883609496e-06 pdrout=1.422132201e-12 pscbe1=9.076987973e+08 lpscbe1=-2.097567017e+01 wpscbe1=-1.361907517e+02 ppscbe1=2.456758588e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=4.442926205e-05 lalpha0=-8.009227281e-12 walpha0=-5.203747270e-11 palpha0=9.387091738e-18 alpha1=0.85 beta0=8.096919820e+01 lbeta0=-1.212820255e-05 wbeta0=-7.664373574e-05 pbeta0=1.384985442e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.651518361e-01 lkt1=2.601077601e-08 wkt1=8.509168044e-08 pkt1=-1.534977333e-14 kt2=1.305987537e-01 lkt2=-2.876834047e-08 wkt2=-1.867869718e-07 pkt2=3.369468862e-14 at=-2.791662271e+05 lat=7.137352880e-02 wat=3.243901624e-01 pat=-7.452659063e-8 ute=1.275482971e+01 lute=-2.538800008e-06 wute=-1.648391105e-05 pute=2.973549199e-12 ua1=3.266627351e-08 lua1=-5.897003590e-15 wua1=-3.828804252e-14 pua1=6.906818278e-21 ub1=-2.845578361e-17 lub1=5.260839563e-24 wub1=3.415755914e-23 pub1=-6.161716251e-30 uc1=-1.159520343e-09 luc1=2.357181089e-16 wuc1=1.530469643e-15 puc1=-2.760829494e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.53 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.023242460e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.610552483e-8 k1=0.90707349 k2=-1.513956257e-01 wk2=4.690385814e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=1.309869106e+00 wnfactor=8.222916387e-7 eta0=0.00069413878 etab=-0.043998 u0=3.195294710e-02 wu0=-5.183386631e-9 ua=-8.937530438e-10 wua=-3.076617972e-16 ub=8.384280427e-19 wub=1.395267750e-24 uc=1.767920239e-11 wuc=7.418974496e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.408109098e+05 wvsat=8.159585085e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=0.0 dwg=0.0 dwb=0.0 pclm=0.14094 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.373633986e+01 wbeta0=1.331235330e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=1.164939156e+05 wat=-8.874902203e-2 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.54 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.945775258e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.361236227e-06 wvth0=-2.039245633e-07 pvth0=4.078571001e-12 k1=4.984927442e-01 lk1=-4.995450494e-07 wk1=8.487159698e-08 pk1=-1.697465124e-12 k2=-3.090125468e-02 lk2=6.522807835e-07 wk2=-9.668171503e-09 pk2=1.933672103e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.324895076e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.633754886e-07 wvoff=-1.297972321e-08 pvoff=2.595995392e-13 nfactor=-3.330107559e+00 lnfactor=1.295906846e-04 wnfactor=6.692877432e-06 pnfactor=-1.338601656e-10 eta0=0.08 etab=-0.07 u0=7.202624000e-02 lu0=-8.963323230e-07 wu0=-4.764111611e-08 pu0=9.528409500e-13 ua=7.842516285e-10 lua=-2.885507167e-14 wua=-1.756257629e-15 pua=3.512583928e-20 ub=2.193434925e-18 lub=-1.969528354e-23 wub=-7.818405599e-25 pub=1.563711690e-29 uc=1.805529429e-10 luc=-3.095139367e-15 wuc=-1.151184154e-16 puc=2.302413320e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.909668800e+00 la0=-1.042135972e-05 wa0=-5.044377618e-07 pa0=1.008895247e-11 ags=5.487759153e-01 lags=-4.295842287e-06 wags=-1.833171611e-07 pags=3.666414900e-12 a1=0.0 a2=0.42385546 b0=-7.783263784e-11 lb0=1.556683189e-15 wb0=9.116085441e-17 pb0=-1.823252732e-21 b1=-4.590399523e-08 lb1=9.180978531e-13 wb1=5.376468719e-14 pb1=-1.075314766e-18 keta=-1.155764801e-02 lketa=2.004897258e-07 wketa=5.702299758e-09 pketa=-1.140482248e-13 dwg=0.0 dwb=0.0 pclm=3.755501550e-01 lpclm=-5.840497280e-06 wpclm=-3.420250992e-07 ppclm=6.840635715e-12 pdiblc1=0.39 pdiblc2=8.871738797e-03 lpdiblc2=-1.144295590e-07 wpdiblc2=-7.708135344e-09 ppdiblc2=1.541657208e-13 pdiblcb=-1.347872257e+01 lpdiblcb=2.252078302e-04 wpdiblcb=1.275932083e-05 ppdiblcb=-2.551914055e-10 drout=0.56 pscbe1=3.292177403e+09 lpscbe1=-5.061426154e+04 wpscbe1=-2.917166737e+03 ppscbe1=5.834447536e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.535595256e-01 lkt1=3.221653494e-06 wkt1=1.537306765e-07 pkt1=-3.074673638e-12 kt2=-9.674096409e-02 lkt2=1.522115958e-06 wkt2=5.923316341e-08 pkt2=-1.184686428e-12 at=-1.333458992e+04 lat=3.066751752e+00 wat=1.795919118e-01 pat=-3.591908456e-6 ute=-4.872681449e+00 lute=7.170103071e-05 wute=3.463045179e-06 pute=-6.926225762e-11 ua1=-3.386311461e-09 lua1=9.480008253e-14 wua1=4.054261752e-15 pua1=-8.108682026e-20 ub1=3.362879455e-19 lub1=-2.556745874e-23 wub1=-7.404831082e-25 pub1=1.480995169e-29 uc1=-5.664850473e-11 luc1=6.448162405e-16 wuc1=9.570211812e-17 puc1=-1.914079782e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.55 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.526519+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.47351598 k2=0.0017121469 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.11141737+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.1493 eta0=0.08 etab=-0.07 u0=0.0272105 ua=-6.5847375e-10 ub=1.20869e-18 uc=2.5799e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.388611 ags=0.333988 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.0015333577 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0031503727 pdiblcb=-2.2185512 drout=0.56 pscbe1=761513800.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.29248 kt2=-0.020636654 at=140000.0 ute=-1.2877 ua1=1.3536e-9 ub1=-9.4206e-19 uc1=-2.4408323e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.56 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.180269700e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.793956050e-8 k1=4.567771039e-01 lk1=1.339175534e-7 k2=1.075904405e-02 lk2=-7.237871452e-08 wk2=1.734723476e-24 pk2=-2.081668171e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.168250686e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.326370282e-8 nfactor=3.356720273e+00 lnfactor=-1.659443288e-6 eta0=0.08 etab=-0.07 u0=2.771774958e-02 lu0=-4.058194965e-9 ua=-6.204091395e-10 lua=-3.045317669e-16 ub=1.202169363e-18 lub=5.216764821e-26 uc=2.622104125e-11 luc=-3.376495022e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.508158685e+00 la0=-9.564282203e-7 ags=3.467182443e-01 lags=-1.018469316e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.282789153e-02 lketa=9.036068682e-08 wketa=3.469446952e-24 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=-3.661419512e-01 lpclm=3.597559432e-06 wpclm=-1.110223025e-22 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=2.956084710e-03 lpdiblc2=1.554379885e-9 pdiblcb=-4.412316820e+00 lpdiblcb=1.755098272e-5 drout=0.56 pscbe1=7.778006919e+08 lpscbe1=-1.303015033e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912498798e-01 lkt1=-9.841442837e-9 kt2=-2.057492397e-02 lkt2=-4.938644046e-10 at=140000.0 ute=-1.489919765e+00 lute=1.617837188e-6 ua1=1.251690039e-09 lua1=8.153195326e-16 ub1=-9.358493930e-19 lub1=-4.968728457e-26 uc1=-3.053243357e-11 luc1=4.899527911e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.57 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.093576859e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.026200865e-7 k1=4.410746075e-01 lk1=1.967336790e-7 k2=1.823098495e-02 lk2=-1.022693997e-07 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.616831167e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.937531150e-8 nfactor=3.523938366e+00 lnfactor=-2.328381042e-6 eta0=0.08 etab=-0.07 u0=2.861607387e-02 lu0=-7.651843391e-9 ua=-2.417916951e-10 lua=-1.819149584e-15 ub=6.901543717e-19 lub=2.100427810e-24 uc=-3.345614174e-12 luc=1.149016872e-16 puc=5.169878828e-38 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.509898072e+00 la0=-9.633864487e-7 ags=1.372902411e-01 lags=7.359469672e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.836687852e-02 lketa=-7.443450054e-08 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=5.092253217e-01 lpclm=9.574807172e-8 pdiblc1=0.39 pdiblc2=1.391985430e-03 lpdiblc2=7.811388567e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.904462922e+08 lpscbe1=2.191502512e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.957403969e-01 lkt1=8.122381345e-9 kt2=-2.369856042e-02 lkt2=1.200190276e-8 at=1.688056304e+05 lat=-1.152337846e-1 ute=-1.748659622e+00 lute=2.652897785e-6 ua1=-7.001213416e-10 lua1=8.623328214e-15 ub1=8.400095403e-19 lub1=-7.153817379e-24 uc1=-6.347849780e-12 luc1=-4.775251223e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.58 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.315090073e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.830878251e-8 k1=5.996005205e-01 lk1=-1.203801308e-7 k2=-5.100121726e-02 lk2=3.622207456e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.003464527e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.101348577e-8 nfactor=2.805264840e+00 lnfactor=-8.907529884e-7 eta0=1.574989903e-01 leta0=-1.550282826e-7 etab=-5.561937938e-02 letab=-2.876686407e-8 u0=2.729087711e-02 lu0=-5.000931709e-9 ua=-9.187605561e-10 lua=-4.649471672e-16 ub=1.549390537e-18 lub=3.816195178e-25 uc=3.803772445e-11 luc=3.211882910e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.999609000e+04 lvsat=2.001173153e-2 a0=1.389139033e+00 la0=-7.218211551e-7 ags=3.400050372e-01 lags=3.304381136e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.723298203e-02 lketa=3.678696011e-8 dwg=0.0 dwb=0.0 pclm=4.258186930e-01 lpclm=2.625939411e-7 pdiblc1=4.413154365e-01 lpdiblc1=-1.026509373e-7 pdiblc2=4.786954283e-03 lpdiblc2=1.020123430e-9 pdiblcb=-6.179303369e-04 lpdiblcb=-4.877367272e-8 drout=7.227638058e-01 ldrout=-3.255912522e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.120046920e-08 lalpha0=-2.401407783e-15 alpha1=1.003059823e+00 lalpha1=-3.061794924e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.267337006e-01 lkt1=7.012110728e-8 kt2=8.365024636e-04 lkt2=-3.707781622e-8 at=1.366949646e+05 lat=-5.099989780e-2 ute=2.021041130e-01 lute=-1.249392435e-06 pute=4.440892099e-28 ua1=5.976024480e-09 lua1=-4.731573803e-15 pua1=3.308722450e-36 ub1=-4.705449676e-18 lub1=3.939269328e-24 uc1=-7.850456210e-11 luc1=9.658912569e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.59 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.922595758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.465539441e-9 k1=3.949806592e-01 lk1=8.431973689e-8 k2=6.610528715e-03 lk2=-2.141219761e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.066022556e-01 ldsub=5.341862293e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.572447639e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.907072680e-9 nfactor=7.446199874e-01 lnfactor=1.170697576e-6 eta0=-4.853186005e-01 leta0=4.880406498e-07 weta0=6.245004514e-23 peta0=1.214306433e-28 etab=-1.685032369e-01 letab=8.416113102e-8 u0=2.366076962e-02 lu0=-1.369404848e-9 ua=-1.285195366e-09 lua=-9.836908175e-17 ub=2.039506695e-18 lub=-1.086882751e-25 uc=6.274221633e-11 luc=7.404677769e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.282663926e+04 lvsat=4.719180553e-2 a0=-1.654509368e-01 la0=8.333766597e-7 ags=2.450957391e-01 lags=4.253845212e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.075565077e-02 lketa=-4.123216624e-08 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=8.767672584e-01 lpclm=-1.885309452e-7 pdiblc1=5.354439199e-01 lpdiblc1=-1.968162250e-7 pdiblc2=1.001082697e-02 lpdiblc2=-4.205791797e-09 ppdiblc2=-3.469446952e-30 pdiblcb=-7.376413933e-02 lpdiblcb=2.440113644e-8 drout=-2.058716915e-01 ldrout=6.034073416e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.759906160e-08 lalpha0=1.201407967e-15 alpha1=5.438803540e-01 lalpha1=1.531795158e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.425064662e-01 lkt1=-1.413906000e-8 kt2=-3.610332050e-02 lkt2=-1.235497918e-10 at=1.213274392e+05 lat=-3.562636363e-2 ute=-8.675146084e-01 lute=-1.793554922e-7 ua1=1.399105300e-09 lua1=-1.528650472e-16 ub1=-8.557691006e-19 lub1=8.808352779e-26 uc1=-3.124743219e-12 luc1=2.117983330e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.60 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.233676712e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.803175043e-8 k1=2.193658629e-01 lk1=1.721958005e-7 k2=7.299517597e-02 lk2=-5.463047764e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.678548315e-01 ldsub=7.280748522e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236272e-03 lcdscd=-1.677929251e-9 cit=0.0 voff='-1.123480252e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.655885130e-8 nfactor=4.230541301e+00 lnfactor=-5.736260754e-07 wnfactor=-3.552713679e-21 eta0=9.800711344e-01 leta0=-2.452271850e-7 etab=4.344132412e-02 letab=-2.189401981e-08 wetab=-4.336808690e-24 petab=-6.938893904e-30 u0=2.299643607e-02 lu0=-1.036978320e-9 ua=-1.853099437e-09 lua=1.858050045e-16 ub=2.473206428e-18 lub=-3.257077184e-25 uc=6.249650872e-11 luc=7.527627645e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.981901101e+04 lvsat=2.367724563e-2 a0=1.5 ags=9.401578928e-01 lags=7.758167506e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.994006187e-02 lketa=-2.581232290e-8 dwg=0.0 dwb=0.0 pclm=7.618388765e-01 lpclm=-1.310218173e-7 pdiblc1=-7.307008025e-02 lpdiblc1=1.076787041e-7 pdiblc2=-5.205115563e-03 lpdiblc2=3.408128906e-09 wpdiblc2=1.734723476e-24 ppdiblc2=4.336808690e-31 pdiblcb=5.341822458e-02 lpdiblcb=-3.923977382e-8 drout=1.497450137e+00 ldrout=-2.489195716e-7 pscbe1=8.085935393e+08 lpscbe1=-4.300129728e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.841313760e-08 lalpha0=-4.209858337e-15 alpha1=0.85 beta0=1.339928056e+01 lbeta0=2.305398613e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.006108499e-01 lkt1=1.493585068e-8 kt2=-4.383320009e-02 lkt2=3.744412390e-9 at=7.157377409e+04 lat=-1.073007741e-2 ute=-1.132701795e+00 lute=-4.665821077e-8 ua1=2.212823246e-09 lua1=-5.600421836e-16 ub1=-2.069402609e-18 lub1=6.953748126e-25 wub1=-7.703719778e-40 uc1=-6.895148964e-11 luc1=5.411894477e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.61 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='7.003489395e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.730716717e-08 wvth0=-9.379950633e-08 pvth0=2.348655219e-14 k1=0.90707349 k2=-1.161455045e-01 lk2=-7.271353509e-09 wk2=-2.735598549e-08 pk2=6.849692563e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586427305e-01 ldsub=-3.187590249e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.036177350e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483740e-8 nfactor=-8.903409017e+00 lnfactor=2.714996879e-06 wnfactor=1.248153545e-05 pnfactor=-3.125264144e-12 eta0=6.941431440e-04 leta0=-7.872186444e-16 etab=-0.043998 u0=-2.848415268e-02 lu0=1.185329778e-08 wu0=2.926963506e-08 pu0=-7.328853192e-15 ua=-3.817646921e-10 lua=-1.826039736e-16 wua=-7.171478440e-16 pua=1.795673658e-22 ub=-5.372131473e-18 lub=1.638694284e-24 wub=5.077677122e-24 pub=-1.271404652e-30 uc=3.857348891e-10 luc=-7.340835366e-17 wuc=-3.085535131e-16 puc=7.725902270e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.346800369e+04 lvsat=2.777139071e-02 wvsat=5.113644001e-02 pvsat=-1.280410435e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.496641316e-01 lketa=1.418505407e-07 wketa=4.125612661e-07 pketa=-1.033016280e-13 dwg=0.0 dwb=0.0 pclm=3.882845217e-01 lpclm=-3.748716880e-08 wpclm=1.193254124e-07 ppclm=-2.987800933e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-7.591454567e-08 lalpha0=2.441676461e-14 walpha0=8.885934963e-14 palpha0=-2.224958141e-20 alpha1=0.85 beta0=1.760852456e+01 lbeta0=-8.234169531e-07 wbeta0=-2.433053621e-06 pbeta0=6.092147292e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.731382297e-01 lkt1=5.813515382e-08 wkt1=2.115698801e-07 pkt1=-5.297519384e-14 kt2=-0.028878939 at=1.784335196e+05 lat=-3.748679593e-02 wat=-2.115698801e-01 pat=5.297519384e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.62 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.391232047e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.815604351e-09 wvth0=1.001292388e-07 pvth0=-1.149644807e-14 k1=0.90707349 k2=-2.434764013e-01 lk2=1.569799430e-08 wk2=1.125392576e-07 pk2=-1.838615024e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.381418108e+01 lnfactor=-4.990871917e-06 wnfactor=-3.724812373e-05 pnfactor=5.845518806e-12 eta0=0.00069413878 etab=-0.043998 u0=7.709010694e-02 lu0=-7.191348489e-09 wu0=-5.804992401e-08 pu0=8.422809387e-15 ua=-1.159830060e-09 lua=-4.224798385e-17 wua=3.978779279e-18 pua=4.948261310e-23 ub=3.506429030e-18 lub=3.708187630e-26 wub=-1.729607062e-24 pub=-4.343185096e-32 uc=-5.336743627e-10 luc=9.244480068e-17 wuc=7.199581972e-16 puc=-1.082752332e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.200223054e+05 lvsat=1.334313669e-03 wvsat=-1.117986258e-02 pvsat=-1.562804210e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=8.218992781e-01 lketa=-1.236062543e-07 wketa=-9.626429543e-07 pketa=1.447728365e-13 dwg=0.0 dwb=0.0 pclm=1.804738837e-01 wpclm=-4.630374500e-8 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.070244599e-07 lalpha0=-2.662288555e-14 walpha0=-2.073384825e-13 palpha0=3.118184172e-20 alpha1=0.85 beta0=9.002901693e+00 lbeta0=7.289599615e-07 wbeta0=5.677125115e-06 pbeta0=-8.537885232e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=2.005260693e-01 lkt1=-6.338782274e-08 wkt1=-4.936630535e-07 pkt1=7.424248028e-14 kt2=-0.028878939 at=-3.807663223e+05 lat=6.338782274e-02 wat=4.936630535e-01 pat=-7.424248028e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.63 nmos lmin=2.0e-05 lmax=0.0001 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.184567870e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.347946121e-06 wvth0=4.768825094e-08 pvth0=-4.768843740e-12 k1=7.025491661e-01 lk1=-1.345419721e-05 wk1=-1.010731850e-07 pk1=1.010735802e-11 k2=-8.210070699e-02 lk2=4.923455350e-06 wk2=3.698691982e-08 pk2=-3.698706444e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.038076407e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.470216738e-07 wvoff=-3.358201432e-09 pvoff=3.358214563e-13 nfactor=4.827326828e+00 lnfactor=-9.857306820e-05 wnfactor=-7.405193935e-07 pnfactor=7.405222890e-11 eta0=0.08 etab=-0.07 u0=1.273385255e-02 lu0=8.504080704e-07 wu0=6.388597617e-09 pu0=-6.388622596e-13 ua=-1.598141021e-09 lua=5.519928788e-14 wua=4.146786129e-16 pua=-4.146802343e-20 ub=1.454467727e-18 lub=-1.443782914e-23 wub=-1.084626123e-25 pub=1.084630364e-29 uc=8.091235261e-11 luc=-3.237547919e-15 wuc=-2.432172464e-17 puc=2.432181974e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.325564408e+00 la0=3.703573706e-06 wa0=2.782269240e-08 pa0=-2.782280118e-12 ags=3.603885030e-01 lags=-1.550856361e-06 wags=-1.165063879e-08 pags=1.165068434e-12 a1=0.0 a2=0.42385546 b0=4.306200292e-11 lb0=-2.529610183e-15 wb0=-1.900341983e-17 pb0=1.900349413e-21 b1=2.539703178e-08 lb1=-1.491909011e-12 wb1=-1.120780327e-14 pb1=1.120784710e-18 keta=-8.836985344e-03 lketa=4.290402119e-07 wketa=3.223117667e-09 pketa=-3.223130269e-13 dwg=0.0 dwb=0.0 pclm=-7.803270971e-02 lpclm=9.490808080e-06 wpclm=7.129865766e-08 ppclm=-7.129893644e-12 pdiblc1=0.39 pdiblc2=-2.157954133e-03 lpdiblc2=3.118293786e-07 wpdiblc2=2.342584101e-09 ppdiblc2=-2.342593260e-13 pdiblcb=3.098273532e+00 lpdiblcb=-3.123285744e-04 wpdiblcb=-2.346334254e-06 ppdiblcb=2.346343429e-10 drout=0.56 pscbe1=-5.389116656e+08 lpscbe1=7.639146525e+04 wpscbe1=5.738825275e+02 ppscbe1=-5.738847714e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.776945549e-01 lkt1=-8.685479070e-07 wkt1=-6.524871155e-09 pkt1=6.524896667e-13 kt2=-4.216347918e-02 lkt2=1.264559762e-06 wkt2=9.499866904e-09 pkt2=-9.499904049e-13 at=2.248345211e+05 lat=-4.983471597e+00 wat=-3.743778532e-02 pat=3.743793170e-6 ute=-8.700717717e-01 lute=-2.453291875e-05 wute=-1.843008689e-07 pute=1.843015895e-11 ua1=7.898140111e-10 lua1=3.311872839e-14 wua1=2.488008247e-16 pua1=-2.488017975e-20 ub1=-3.896016502e-20 lub1=-5.305119093e-23 wub1=-3.985412695e-25 pub1=3.985428277e-29 uc1=1.167240467e-10 luc1=-8.290600883e-15 wuc1=-6.228223236e-17 puc1=6.228247589e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.64 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='8.754073007e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.791242821e-06 wvth0=-3.179216729e-07 pvth0=2.543497691e-12 k1=-2.659376817e-01 lk1=5.915918420e-06 wk1=6.738212336e-07 pk1=-5.390833333e-12 k2=2.723092720e-01 lk2=-2.164882804e-06 wk2=-2.465794655e-07 pk2=1.972732136e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.359860461e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.965590152e-07 wvoff=2.238800955e-08 pvoff=-1.791128301e-13 nfactor=-2.268356294e+00 lnfactor=4.334336866e-05 wnfactor=4.936795957e-06 pnfactor=-3.949629794e-11 eta0=0.08 etab=-0.07 u0=7.394962174e-02 lu0=-3.739312490e-07 wu0=-4.259065078e-08 pu0=3.407418592e-13 ua=2.375324172e-09 lua=-2.427156959e-14 wua=-2.764524086e-15 pua=2.211727362e-20 ub=4.151751246e-19 lub=6.348429268e-24 wub=7.230840821e-25 pub=-5.784955383e-30 uc=-1.521392765e-10 luc=1.423575786e-15 wuc=1.621448310e-16 puc=-1.297222046e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.592162434e+00 la0=-1.628491062e-06 wa0=-1.854846160e-07 pa0=1.483949452e-12 ags=2.487516684e-01 lags=6.819239801e-07 wags=7.767092527e-08 pags=-6.213977715e-13 a1=0.0 a2=0.42385546 b0=-1.390294406e-10 lb0=1.112289885e-15 wb0=1.266894655e-16 pb0=-1.013565260e-21 b1=-8.199653713e-08 lb1=6.560043577e-13 wb1=7.471868848e-14 pb1=-5.977787229e-19 keta=2.204704258e-02 lketa=-1.886524222e-07 wketa=-2.148745111e-08 pketa=1.719080105e-13 dwg=0.0 dwb=0.0 pclm=6.051535595e-01 lpclm=-4.173184431e-06 wpclm=-4.753243844e-07 ppclm=3.802780927e-12 pdiblc1=0.39 pdiblc2=2.028876990e-02 lpdiblc2=-1.371138787e-07 wpdiblc2=-1.561722734e-08 ppdiblc2=1.249439250e-13 pdiblcb=-1.938438460e+01 lpdiblcb=1.373333791e-04 wpdiblcb=1.564222836e-05 ppdiblcb=-1.251439430e-10 drout=0.56 pscbe1=4.960051090e+09 lpscbe1=-3.358993994e+04 wpscbe1=-3.825883517e+03 ppscbe1=3.060856406e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.402161020e-01 lkt1=3.819074806e-07 wkt1=4.349914103e-08 pkt1=-3.480101364e-13 kt2=4.886458281e-02 lkt2=-5.560370694e-07 wkt2=-6.333244603e-08 pkt2=5.066843312e-13 at=-1.338956671e+05 lat=2.191272430e+00 wat=2.495852354e-01 pat=-1.996779471e-6 ute=-2.636049241e+00 lute=1.078732113e-05 wute=1.228672459e-06 pute=-9.829860083e-12 ua1=3.173832347e-09 lua1=-1.456257049e-14 wua1=-1.658672165e-15 pua1=1.327002586e-20 ub1=-3.857796760e-18 lub1=2.332703413e-23 wub1=2.656941796e-24 pub1=-2.125657324e-29 uc1=-4.800665152e-10 luc1=3.645443700e-15 wuc1=4.152148824e-16 puc1=-3.321881408e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.65 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.180269700e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.793956050e-8 k1=4.567771039e-01 lk1=1.339175534e-7 k2=1.075904405e-02 lk2=-7.237871452e-08 pk2=1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.168250686e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.326370282e-8 nfactor=3.356720273e+00 lnfactor=-1.659443288e-6 eta0=0.08 etab=-0.07 u0=2.771774958e-02 lu0=-4.058194965e-9 ua=-6.204091395e-10 lua=-3.045317669e-16 ub=1.202169363e-18 lub=5.216764821e-26 uc=2.622104125e-11 luc=-3.376495022e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.508158685e+00 la0=-9.564282203e-7 ags=3.467182443e-01 lags=-1.018469316e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.282789153e-02 lketa=9.036068682e-08 wketa=3.469446952e-24 pketa=-2.081668171e-29 dwg=0.0 dwb=0.0 pclm=-3.661419512e-01 lpclm=3.597559432e-06 wpclm=-1.110223025e-22 pdiblc1=0.39 pdiblc2=2.956084710e-03 lpdiblc2=1.554379885e-9 pdiblcb=-4.412316820e+00 lpdiblcb=1.755098272e-5 drout=0.56 pscbe1=7.778006919e+08 lpscbe1=-1.303015033e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912498798e-01 lkt1=-9.841442837e-9 kt2=-2.057492397e-02 lkt2=-4.938644046e-10 at=140000.0 ute=-1.489919765e+00 lute=1.617837188e-6 ua1=1.251690039e-09 lua1=8.153195326e-16 ub1=-9.358493930e-19 lub1=-4.968728457e-26 uc1=-3.053243357e-11 luc1=4.899527911e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.66 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.093576859e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.026200865e-7 k1=4.410746075e-01 lk1=1.967336790e-7 k2=1.823098495e-02 lk2=-1.022693997e-07 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.616831167e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.937531150e-8 nfactor=3.523938366e+00 lnfactor=-2.328381042e-6 eta0=0.08 etab=-0.07 u0=2.861607387e-02 lu0=-7.651843391e-9 ua=-2.417916951e-10 lua=-1.819149584e-15 ub=6.901543717e-19 lub=2.100427810e-24 uc=-3.345614173e-12 luc=1.149016872e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.509898072e+00 la0=-9.633864487e-7 ags=1.372902411e-01 lags=7.359469672e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.836687852e-02 lketa=-7.443450054e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.092253217e-01 lpclm=9.574807172e-8 pdiblc1=0.39 pdiblc2=1.391985430e-03 lpdiblc2=7.811388567e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.904462922e+08 lpscbe1=2.191502512e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.957403969e-01 lkt1=8.122381345e-9 kt2=-2.369856042e-02 lkt2=1.200190276e-8 at=1.688056304e+05 lat=-1.152337846e-1 ute=-1.748659622e+00 lute=2.652897785e-6 ua1=-7.001213416e-10 lua1=8.623328214e-15 ub1=8.400095403e-19 lub1=-7.153817379e-24 uc1=-6.347849780e-12 luc1=-4.775251223e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.67 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.315090073e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.830878251e-8 k1=5.996005205e-01 lk1=-1.203801308e-7 k2=-5.100121726e-02 lk2=3.622207456e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.003464527e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.101348577e-8 nfactor=2.805264840e+00 lnfactor=-8.907529884e-7 eta0=1.574989903e-01 leta0=-1.550282826e-07 weta0=-1.110223025e-22 etab=-5.561937937e-02 letab=-2.876686407e-8 u0=2.729087711e-02 lu0=-5.000931709e-9 ua=-9.187605561e-10 lua=-4.649471672e-16 ub=1.549390537e-18 lub=3.816195178e-25 uc=3.803772445e-11 luc=3.211882910e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.999609000e+04 lvsat=2.001173153e-2 a0=1.389139033e+00 la0=-7.218211551e-7 ags=3.400050372e-01 lags=3.304381136e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.723298203e-02 lketa=3.678696011e-08 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=4.258186930e-01 lpclm=2.625939411e-7 pdiblc1=4.413154365e-01 lpdiblc1=-1.026509373e-7 pdiblc2=4.786954283e-03 lpdiblc2=1.020123430e-9 pdiblcb=-6.179303369e-04 lpdiblcb=-4.877367272e-8 drout=7.227638058e-01 ldrout=-3.255912522e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.120046920e-08 lalpha0=-2.401407783e-15 alpha1=1.003059823e+00 lalpha1=-3.061794924e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.267337006e-01 lkt1=7.012110728e-8 kt2=8.365024636e-04 lkt2=-3.707781622e-8 at=1.366949646e+05 lat=-5.099989780e-2 ute=2.021041130e-01 lute=-1.249392435e-6 ua1=5.976024480e-09 lua1=-4.731573803e-15 ub1=-4.705449676e-18 lub1=3.939269328e-24 uc1=-7.850456210e-11 luc1=9.658912569e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.68 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.922595758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.465539441e-9 k1=3.949806592e-01 lk1=8.431973689e-8 k2=6.610528715e-03 lk2=-2.141219761e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.066022556e-01 ldsub=5.341862293e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.572447639e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.907072680e-9 nfactor=7.446199874e-01 lnfactor=1.170697576e-6 eta0=-4.853186005e-01 leta0=4.880406498e-07 weta0=-1.179611964e-22 peta0=-2.255140519e-29 etab=-1.685032369e-01 letab=8.416113102e-8 u0=2.366076962e-02 lu0=-1.369404848e-9 ua=-1.285195366e-09 lua=-9.836908175e-17 ub=2.039506695e-18 lub=-1.086882751e-25 uc=6.274221633e-11 luc=7.404677769e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.282663926e+04 lvsat=4.719180553e-2 a0=-1.654509368e-01 la0=8.333766597e-7 ags=2.450957391e-01 lags=4.253845212e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.075565077e-02 lketa=-4.123216624e-08 wketa=1.387778781e-23 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=8.767672584e-01 lpclm=-1.885309452e-7 pdiblc1=5.354439199e-01 lpdiblc1=-1.968162250e-7 pdiblc2=1.001082697e-02 lpdiblc2=-4.205791797e-9 pdiblcb=-7.376413933e-02 lpdiblcb=2.440113644e-8 drout=-2.058716915e-01 ldrout=6.034073416e-07 pdrout=2.220446049e-28 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.759906160e-08 lalpha0=1.201407967e-15 alpha1=5.438803540e-01 lalpha1=1.531795158e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.425064662e-01 lkt1=-1.413906000e-8 kt2=-3.610332050e-02 lkt2=-1.235497918e-10 at=1.213274392e+05 lat=-3.562636363e-2 ute=-8.675146084e-01 lute=-1.793554922e-7 ua1=1.399105300e-09 lua1=-1.528650472e-16 ub1=-8.557691006e-19 lub1=8.808352779e-26 uc1=-3.124743219e-12 luc1=2.117983330e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.69 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.233676712e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.803175043e-8 k1=2.193658629e-01 lk1=1.721958005e-7 k2=7.299517597e-02 lk2=-5.463047764e-08 pk2=-1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.678548315e-01 ldsub=7.280748522e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236272e-03 lcdscd=-1.677929251e-9 cit=0.0 voff='-1.123480252e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.655885130e-8 nfactor=4.230541301e+00 lnfactor=-5.736260754e-7 eta0=9.800711344e-01 leta0=-2.452271850e-7 etab=4.344132412e-02 letab=-2.189401981e-08 wetab=-1.040834086e-23 petab=4.553649124e-30 u0=2.299643607e-02 lu0=-1.036978320e-9 ua=-1.853099437e-09 lua=1.858050045e-16 ub=2.473206428e-18 lub=-3.257077184e-25 uc=6.249650872e-11 luc=7.527627645e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.981901101e+04 lvsat=2.367724563e-2 a0=1.5 ags=9.401578928e-01 lags=7.758167506e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.994006187e-02 lketa=-2.581232290e-8 dwg=0.0 dwb=0.0 pclm=7.618388765e-01 lpclm=-1.310218173e-7 pdiblc1=-7.307008025e-02 lpdiblc1=1.076787041e-7 pdiblc2=-5.205115563e-03 lpdiblc2=3.408128906e-09 ppdiblc2=4.336808690e-31 pdiblcb=5.341822458e-02 lpdiblcb=-3.923977382e-8 drout=1.497450137e+00 ldrout=-2.489195716e-7 pscbe1=8.085935393e+08 lpscbe1=-4.300129728e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.841313760e-08 lalpha0=-4.209858337e-15 alpha1=0.85 beta0=1.339928056e+01 lbeta0=2.305398613e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.006108499e-01 lkt1=1.493585068e-8 kt2=-4.383320009e-02 lkt2=3.744412390e-9 at=7.157377409e+04 lat=-1.073007741e-2 ute=-1.132701795e+00 lute=-4.665821077e-8 ua1=2.212823246e-09 lua1=-5.600421836e-16 ub1=-2.069402609e-18 lub1=6.953748126e-25 pub1=1.925929944e-46 uc1=-6.895148964e-11 luc1=5.411894477e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.70 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.974130494e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.153294672e-8 k1=0.90707349 k2=-1.461660539e-01 lk2=2.455218805e-10 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586427305e-01 ldsub=-3.187590249e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.036177350e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483740e-8 nfactor=4.793869483e+00 lnfactor=-7.146783822e-07 wnfactor=3.552713679e-21 eta0=6.941431440e-04 leta0=-7.872186444e-16 etab=-0.043998 u0=3.636442136e-03 lu0=3.810589922e-9 ua=-1.168765120e-09 lua=1.445385052e-17 ub=2.001282801e-19 lub=2.434505921e-25 uc=4.712723814e-11 luc=1.137595467e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.295853029e+05 lvsat=1.372012403e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.969180267e-01 lketa=2.848699075e-8 dwg=0.0 dwb=0.0 pclm=5.192326259e-01 lpclm=-7.027539555e-8 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.16e-8 alpha1=0.85 beta0=1.493848343e+01 lbeta0=-1.548626842e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.24096074 kt2=-0.028878939 at=-5.374397014e+04 lat=2.064835789e-2 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.71 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.638575314e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.479833270e-09 wvth0=-1.353391853e-08 pvth0=2.441397097e-15 k1=0.90707349 k2=9.928057558e-03 lk2=-2.791245099e-08 wk2=-1.183735283e-07 pk2=2.135351914e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587413353e-01 ldsub=-2.097501524e-11 wdsub=-1.059549248e-10 pdsub=1.911331483e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-1.099938796e+01 lnfactor=2.134283121e-06 wnfactor=3.587882554e-06 pnfactor=-6.472217217e-13 eta0=-1.564415634e-02 leta0=2.947281677e-09 weta0=1.488814215e-08 peta0=-2.685686850e-15 etab=-0.043998 u0=4.168639461e-03 lu0=3.714586315e-09 wu0=8.399179866e-09 pu0=-1.515136455e-15 ua=-3.916177980e-09 lua=5.100624037e-16 wua=2.515678770e-15 pua=-4.538058091e-22 ub=1.563199941e-17 lub=-2.540320073e-24 wub=-1.277893607e-23 pub=2.305205056e-30 uc=1.618364514e-10 luc=-9.316555023e-18 wuc=8.617953193e-17 puc=-1.554601194e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.230348001e+05 lvsat=-1.294110242e-01 wvsat=-6.517943742e-01 pvsat=1.175778390e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.700210004e-01 lketa=1.499087093e-07 wketa=5.791058641e-07 pketa=-1.044654859e-13 dwg=0.0 dwb=0.0 pclm=9.247073827e-02 lpclm=6.708608112e-09 wpclm=3.388841723e-08 ppclm=-6.113165473e-15 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.050948000e-08 lalpha0=7.596171207e-15 alpha1=0.85 beta0=1.994049915e+01 lbeta0=-1.057181302e-06 wbeta0=-4.289673068e-06 pbeta0=7.738184143e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-8.119715551e-01 lkt1=1.030052119e-07 wkt1=4.289673068e-07 pkt1=-7.738184143e-14 kt2=-0.028878939 at=4.669687501e+05 lat=-7.328353044e-02 wat=-2.788287494e-01 pat=5.029819693e-8 ute=-1.421678289e-01 lute=-2.122977251e-07 wute=-1.072418267e-06 pute=1.934546036e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.72 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.73 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.522125473e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.944806751e-7 k1=6.310052922e-01 lk1=-1.259976076e-6 k2=-5.591980128e-02 lk2=4.610781196e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.061847177e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.186326434e-8 nfactor=4.303155891e+00 lnfactor=-9.231298284e-6 eta0=0.08 etab=-0.07 u0=1.725597206e-02 lu0=7.964011574e-8 ua=-1.304613965e-09 lua=5.169374362e-15 ub=1.377693304e-18 lub=-1.352092512e-24 uc=6.369640755e-11 luc=-3.031940783e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.345258486e+00 la0=3.468370644e-7 ags=3.521416882e-01 lags=-1.452366039e-7 a1=0.0 a2=0.42385546 b0=2.961057888e-11 lb0=-2.368962087e-16 b1=1.746367474e-08 lb1=-1.397162262e-13 keta=-6.555526381e-03 lketa=4.017931312e-8 dwg=0.0 dwb=0.0 pclm=-2.756450521e-02 lpclm=8.888074800e-07 ppclm=2.220446049e-28 pdiblc1=0.39 pdiblc2=-4.997740590e-04 lpdiblc2=2.920260128e-8 pdiblcb=1.437438940e+00 lpdiblcb=-2.924935061e-05 wpdiblcb=-8.326672685e-23 ppdiblcb=-1.243449788e-26 drout=0.56 pscbe1=-1.326933481e+08 lpscbe1=7.154006820e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.823131346e-01 lkt1=-8.133889864e-8 kt2=-3.543907171e-02 lkt2=1.184251295e-7 at=1.983344738e+05 lat=-4.666985988e-1 ute=-1.000527719e+00 lute=-2.297490531e-6 ua1=9.659257545e-10 lua1=3.101545545e-15 ub1=-3.210645264e-19 lub1=-4.968206598e-24 uc1=7.263804922e-11 luc1=-7.764089229e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.74 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.180269700e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.793956050e-8 k1=4.567771039e-01 lk1=1.339175534e-7 k2=1.075904405e-02 lk2=-7.237871452e-08 wk2=-3.469446952e-24 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.168250686e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.326370282e-8 nfactor=3.356720273e+00 lnfactor=-1.659443288e-06 wnfactor=3.552713679e-21 eta0=0.08 etab=-0.07 u0=2.771774958e-02 lu0=-4.058194965e-9 ua=-6.204091395e-10 lua=-3.045317669e-16 ub=1.202169363e-18 lub=5.216764821e-26 uc=2.622104125e-11 luc=-3.376495022e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.508158685e+00 la0=-9.564282203e-7 ags=3.467182443e-01 lags=-1.018469316e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.282789153e-02 lketa=9.036068682e-08 wketa=-3.469446952e-24 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=-3.661419512e-01 lpclm=3.597559432e-06 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=2.956084710e-03 lpdiblc2=1.554379885e-9 pdiblcb=-4.412316820e+00 lpdiblcb=1.755098272e-5 drout=0.56 pscbe1=7.778006919e+08 lpscbe1=-1.303015033e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912498798e-01 lkt1=-9.841442837e-9 kt2=-2.057492397e-02 lkt2=-4.938644046e-10 at=140000.0 ute=-1.489919765e+00 lute=1.617837188e-6 ua1=1.251690039e-09 lua1=8.153195326e-16 ub1=-9.358493930e-19 lub1=-4.968728457e-26 uc1=-3.053243357e-11 luc1=4.899527911e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.75 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.093576859e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.026200865e-7 k1=4.410746075e-01 lk1=1.967336790e-7 k2=1.823098495e-02 lk2=-1.022693997e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.616831167e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.937531150e-8 nfactor=3.523938366e+00 lnfactor=-2.328381042e-6 eta0=0.08 etab=-0.07 u0=2.861607387e-02 lu0=-7.651843391e-9 ua=-2.417916951e-10 lua=-1.819149584e-15 ub=6.901543717e-19 lub=2.100427810e-24 uc=-3.345614173e-12 luc=1.149016872e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.509898072e+00 la0=-9.633864487e-7 ags=1.372902411e-01 lags=7.359469672e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.836687852e-02 lketa=-7.443450054e-08 wketa=1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.092253217e-01 lpclm=9.574807172e-8 pdiblc1=0.39 pdiblc2=1.391985430e-03 lpdiblc2=7.811388567e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.904462922e+08 lpscbe1=2.191502512e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.957403969e-01 lkt1=8.122381345e-9 kt2=-2.369856042e-02 lkt2=1.200190276e-8 at=1.688056304e+05 lat=-1.152337846e-1 ute=-1.748659622e+00 lute=2.652897785e-6 ua1=-7.001213416e-10 lua1=8.623328214e-15 pua1=-3.308722450e-36 ub1=8.400095403e-19 lub1=-7.153817379e-24 pub1=-3.081487911e-45 uc1=-6.347849780e-12 luc1=-4.775251223e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.76 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.315090073e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.830878251e-8 k1=5.996005205e-01 lk1=-1.203801308e-7 k2=-5.100121726e-02 lk2=3.622207456e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.003464527e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.101348577e-8 nfactor=2.805264840e+00 lnfactor=-8.907529884e-7 eta0=1.574989903e-01 leta0=-1.550282826e-7 etab=-5.561937937e-02 letab=-2.876686407e-8 u0=2.729087711e-02 lu0=-5.000931709e-09 wu0=2.775557562e-23 ua=-9.187605561e-10 lua=-4.649471672e-16 ub=1.549390537e-18 lub=3.816195178e-25 uc=3.803772445e-11 luc=3.211882910e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.999609000e+04 lvsat=2.001173153e-2 a0=1.389139033e+00 la0=-7.218211551e-7 ags=3.400050372e-01 lags=3.304381136e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.723298203e-02 lketa=3.678696011e-8 dwg=0.0 dwb=0.0 pclm=4.258186930e-01 lpclm=2.625939411e-7 pdiblc1=4.413154365e-01 lpdiblc1=-1.026509373e-07 wpdiblc1=-4.440892099e-22 pdiblc2=4.786954283e-03 lpdiblc2=1.020123430e-9 pdiblcb=-6.179303369e-04 lpdiblcb=-4.877367272e-8 drout=7.227638058e-01 ldrout=-3.255912522e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.120046920e-08 lalpha0=-2.401407783e-15 alpha1=1.003059823e+00 lalpha1=-3.061794924e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.267337006e-01 lkt1=7.012110728e-8 kt2=8.365024636e-04 lkt2=-3.707781622e-8 at=1.366949646e+05 lat=-5.099989780e-2 ute=2.021041130e-01 lute=-1.249392435e-6 ua1=5.976024480e-09 lua1=-4.731573803e-15 ub1=-4.705449676e-18 lub1=3.939269328e-24 uc1=-7.850456210e-11 luc1=9.658912569e-17 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.77 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.921197749e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.325683854e-09 wvth0=1.050243264e-10 pvth0=-1.050653909e-16 k1=-1.818473065e-01 lk1=6.613732423e-07 wk1=4.333373946e-07 pk1=-4.335068295e-13 k2=1.824172536e-01 lk2=-1.972876630e-07 wk2=-1.320733957e-07 pk2=1.321250364e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.867310762e-01 ldsub=7.329757195e-08 wdsub=1.492806455e-08 pdsub=-1.493390142e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.454909514e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.851335601e-09 wvoff=-8.829957640e-09 pvoff=8.833410154e-15 nfactor=4.896190415e-01 lnfactor=1.425798228e-06 wnfactor=1.915674206e-07 pnfactor=-1.916423235e-13 eta0=-4.853186004e-01 leta0=4.880406497e-07 weta0=-9.826697095e-17 peta0=9.830592243e-23 etab=-1.705399596e-01 letab=8.619865007e-08 wetab=1.530071632e-09 petab=-1.530669890e-15 u0=1.419538590e-02 lu0=8.099679840e-09 wu0=7.110793798e-09 pu0=-7.113574119e-15 ua=-1.039313727e-09 lua=-3.443468605e-16 wua=-1.847166143e-16 pua=1.847888385e-22 ub=4.789547535e-19 lub=1.452473842e-24 wub=1.172352161e-24 pub=-1.172810551e-30 uc=-1.002151541e-10 luc=1.704257645e-16 wuc=1.224204208e-16 puc=-1.224682872e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.012648825e+06 lvsat=-9.230095803e-01 wvsat=-7.285711582e-01 pvsat=7.288560295e-7 a0=-9.175719024e-01 la0=1.585791705e-06 wa0=5.650248584e-07 pa0=-5.652457832e-13 ags=-5.874522816e+00 lags=6.547395847e-06 wags=4.597314483e-06 pags=-4.599112032e-12 a1=0.0 a2=0.42385546 b0=-1.499134706e-16 lb0=1.499720867e-22 wb0=1.126212954e-22 pb0=-1.126653304e-28 b1=3.345420305e-17 lb1=-3.346728365e-23 wb1=-2.513220241e-23 pb1=2.514202910e-29 keta=2.106363115e-01 lketa=-2.011753403e-07 wketa=-1.201090673e-07 pketa=1.201560300e-13 dwg=0.0 dwb=0.0 pclm=5.626883191e-01 lpclm=1.256707989e-07 wpclm=2.359492905e-07 ppclm=-2.360415467e-13 pdiblc1=-1.755336640e-01 lpdiblc1=5.144393512e-07 wpdiblc1=5.341162221e-07 ppdiblc1=-5.343250616e-13 pdiblc2=-1.524417998e-04 lpdiblc2=5.961450816e-09 wpdiblc2=7.635074361e-09 ppdiblc2=-7.638059675e-15 pdiblcb=-5.274169803e-01 lpdiblcb=4.782313557e-07 wpdiblcb=3.408030676e-07 ppdiblcb=-3.409363216e-13 drout=-2.058723435e-01 ldrout=6.034079938e-07 wdrout=4.897804500e-13 pdrout=-4.899719535e-19 pscbe1=-1.566202475e+09 lpscbe1=2.367127660e+03 wpscbe1=1.777590680e+03 ppscbe1=-1.778285718e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.525037326e-05 lalpha0=-2.523143490e-11 walpha0=-1.894840734e-11 palpha0=1.895581616e-17 alpha1=5.438803540e-01 lalpha1=1.531795158e-7 beta0=4.095981785e+01 lbeta0=-2.711041387e-05 wbeta0=-2.035852136e-05 pbeta0=2.036648154e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.958659293e-01 lkt1=3.924126668e-08 wkt1=4.008586980e-08 pkt1=-4.010154338e-14 kt2=-3.850419620e-02 lkt2=2.278264658e-09 wkt2=1.803638668e-09 pkt2=-1.804343891e-15 at=-1.359522091e+05 lat=2.217538810e-01 wat=1.932792776e-01 pat=-1.933548498e-7 ute=-1.417159919e+00 lute=3.705047297e-07 wute=4.129166424e-07 pute=-4.130780928e-13 ua1=-3.081215028e-10 lua1=1.555029282e-15 wua1=1.282540478e-15 pua1=-1.283041951e-21 ub1=-5.438363797e-19 lub1=-2.239711588e-25 wub1=-2.343369611e-25 pub1=2.344285869e-31 uc1=-2.212098164e-10 luc1=2.393501777e-16 wuc1=1.638346665e-16 puc1=-1.638987259e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.78 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.780327363e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.723343472e-09 wvth0=3.405750721e-08 pvth0=-1.709458225e-14 k1=1.373021793e+00 lk1=-1.166692614e-07 wk1=-8.666747886e-07 pk1=2.170075668e-13 k2=-2.806519574e-01 lk2=3.442800261e-08 wk2=2.656745798e-07 pk2=-6.690447082e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.075971904e-01 ldsub=6.285635619e-08 wdsub=-2.985612920e-08 pdsub=7.475706071e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236264e-03 lcdscd=-1.677929247e-09 wcdscd=6.014522214e-18 pcdscd=-3.009613392e-24 cit=0.0 voff='-1.358556500e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.067275367e-08 wvoff=1.765991510e-08 pvoff=-4.421883755e-15 nfactor=4.740543194e+00 lnfactor=-7.013259600e-07 wnfactor=-3.831348427e-07 pnfactor=9.593351675e-14 eta0=9.800711345e-01 leta0=-2.452271851e-07 weta0=-6.809930397e-17 peta0=8.321032752e-23 etab=4.751476948e-02 letab=-2.291397385e-08 wetab=-3.060143235e-09 petab=7.662323176e-16 u0=5.084947544e-02 lu0=-1.024169668e-08 wu0=-2.092437300e-08 pu0=6.914971032e-15 ua=-2.344862712e-09 lua=3.089381018e-16 wua=3.694332260e-16 pua=-9.250275429e-23 ub=5.594310312e-18 lub=-1.107204041e-24 wub=-2.344704324e-24 pub=5.870928606e-31 uc=3.884112496e-10 luc=-7.407849027e-17 wuc=-2.448408418e-16 puc=6.130594323e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.529631311e+06 lvsat=3.491245192e-01 wvsat=1.216599099e+00 pvsat=-2.444896607e-7 a0=3.004241928e+00 la0=-3.766486400e-07 wa0=-1.130049715e-06 pa0=2.829542776e-13 ags=1.317939500e+01 lags=-2.987013144e-06 wags=-9.194628965e-06 pags=2.302252341e-12 a1=0.0 a2=0.42385546 b0=2.998269411e-16 lb0=-7.507396761e-23 wb0=-2.252425909e-22 pb0=5.639871758e-29 b1=-6.690840611e-17 lb1=1.675326271e-23 wb1=5.026440482e-23 pb1=-1.258575459e-29 keta=-2.998212595e-01 lketa=5.425303410e-08 wketa=2.402181346e-07 pketa=-6.014845893e-14 dwg=0.0 dwb=0.0 pclm=1.389996755e+00 lpclm=-2.883068968e-07 wpclm=-4.718985813e-07 ppclm=1.181591577e-13 pdiblc1=1.348885088e+00 lpdiblc1=-2.483660726e-07 wpdiblc1=-1.068232445e-06 ppdiblc1=2.674757901e-13 pdiblc2=1.512142197e-02 lpdiblc2=-1.681453152e-09 wpdiblc2=-1.527014871e-08 ppdiblc2=3.823507804e-15 pdiblcb=9.607239065e-01 lpdiblcb=-2.664209508e-07 wpdiblcb=-6.816061351e-07 ppdiblcb=1.706680418e-13 drout=1.497451439e+00 ldrout=-2.489198968e-07 wdrout=-9.777256533e-13 pdrout=2.443548919e-19 pscbe1=5.540998489e+09 lpscbe1=-1.189251738e+03 wpscbe1=-3.555181360e+03 ppscbe1=8.901854158e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.040713526e-05 lalpha0=1.262690145e-11 walpha0=3.789681467e-11 palpha0=-9.489021322e-18 alpha1=0.85 beta0=-4.080035513e+01 lbeta0=1.380164084e-05 wbeta0=4.071704272e-05 pbeta0=-1.019518104e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.938919237e-01 lkt1=-1.178560795e-08 wkt1=-8.017173955e-08 pkt1=2.007428202e-14 kt2=-3.903144869e-02 lkt2=2.542097059e-09 wkt2=-3.607277325e-09 pkt2=9.032297739e-16 at=5.861330707e+05 lat=-1.395710943e-01 wat=-3.865585551e-01 pat=9.679078318e-8 ute=-3.341117355e-02 lute=-3.219106888e-07 wute=-8.258332850e-07 pute=2.067812221e-13 ua1=5.627276849e-09 lua1=-1.414990635e-15 wua1=-2.565080954e-15 pua1=6.422731846e-22 ub1=-2.693268055e-18 lub1=8.515851064e-25 wub1=4.686739252e-25 pub1=-1.173517335e-31 uc1=3.672186568e-10 luc1=-5.509413438e-17 wuc1=-3.276693331e-16 puc1=8.204545200e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.79 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='1.107519298e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.278553263e-07 wvth0=-3.832132387e-07 pvth0=8.738625709e-14 k1=9.070734931e-01 lk1=-5.682059268e-16 wk1=-2.366306262e-15 pk1=4.268603249e-22 k2=-9.384767530e-02 lk2=-1.234610839e-08 wk2=-3.930376341e-08 pk2=9.459361507e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587256360e-01 ldsub=-2.394643062e-11 wdsub=-6.228214134e-11 pdsub=1.559491276e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000032e-03 lcdscd=-6.012607079e-18 wcdscd=-2.404461352e-17 pcdscd=4.516923294e-24 cit=0.0 voff='-1.036177363e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483713e-08 wvoff=9.905569698e-16 pvoff=-2.022012557e-22 nfactor=2.841984073e+01 lnfactor=-6.630408950e-06 wnfactor=-1.774882189e-05 pnfactor=4.444145263e-12 eta0=-1.095530700e-02 leta0=2.916916596e-09 weta0=8.751556224e-09 peta0=-2.191310848e-15 etab=-4.399799986e-02 letab=-2.453373615e-17 wetab=-1.021713825e-16 petab=1.843078468e-23 u0=-1.016275855e-02 lu0=5.035217600e-09 wu0=1.036653912e-08 pu0=-9.199917459e-16 ua=-7.974223360e-10 lua=-7.852704133e-17 wua=-2.789682958e-16 pua=6.985115116e-23 ub=1.312346779e-18 lub=-3.503891036e-26 wub=-8.355452494e-25 pub=2.092130108e-31 uc=-5.098201056e-10 luc=1.508305570e-16 wuc=4.184022364e-16 puc=-1.047641543e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.531072018e+05 lvsat=5.453347092e-02 wvsat=3.626188827e-01 pvsat=-3.066070035e-8 a0=1.500000010e+00 la0=-1.735765309e-15 wa0=-7.228631915e-15 pa0=1.303980035e-21 ags=1.250000002e+00 lags=-3.716431607e-16 wags=-1.547714845e-15 pags=2.791940013e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.473165337e-03 lketa=-2.193955123e-08 wketa=-1.512935219e-07 pketa=3.788253625e-14 dwg=0.0 dwb=0.0 pclm=1.352260278e+00 lpclm=-2.788580224e-07 wpclm=-6.258053592e-07 ppclm=1.566960298e-13 pdiblc1=3.569721484e-01 lpdiblc1=2.971594082e-16 wpdiblc1=1.237526526e-15 ppdiblc1=-2.232385388e-22 pdiblc2=8.406112144e-03 lpdiblc2=-7.967522475e-18 wpdiblc2=-3.318090247e-17 ppdiblc2=5.985534984e-24 pdiblcb=-1.032957699e-01 lpdiblcb=-2.359124007e-17 wpdiblcb=-9.824629998e-17 ppdiblcb=1.772271219e-23 drout=5.033266687e-01 ldrout=-1.573879693e-15 wdrout=-6.554454757e-15 pdrout=1.182364873e-21 pscbe1=7.914198809e+08 lpscbe1=-1.554861069e-07 wpscbe1=-6.475257874e-07 ppscbe1=1.168074608e-13 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.625738297e-07 lalpha0=-3.529857855e-14 walpha0=-1.059054618e-13 palpha0=2.651777475e-20 alpha1=0.85 beta0=1.129890585e+01 lbeta0=7.564547859e-07 wbeta0=2.734203540e-06 pbeta0=-6.846199589e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-8.415575641e-02 lkt1=-3.926255663e-08 wkt1=-1.177984895e-07 pkt1=2.949568157e-14 kt2=-2.887893895e-02 lkt2=-9.431011527e-18 wkt2=-3.927569381e-17 pkt2=7.084999254e-24 at=-1.712221660e+05 lat=5.006384084e-02 wat=8.825455484e-02 pat=-2.209814624e-8 ute=-1.263938142e+00 lute=-1.379781053e-08 wute=-4.139723373e-08 pute=1.036549478e-14 ua1=-2.384732614e-11 lua1=-1.779476610e-24 wua1=-7.410666647e-24 pua1=1.336817561e-30 ub1=7.077531840e-19 lub1=-2.527832356e-33 wub1=-1.052720857e-32 pub1=1.899013918e-39 uc1=1.471862498e-10 luc1=3.660129454e-26 wuc1=1.524266394e-25 puc1=-2.749641414e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.80 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='-2.420807557e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.156003771e-07 wvth0=5.919207722e-07 pvth0=-8.851914227e-14 k1=0.90707349 k2=-3.410479518e-01 lk2=3.224659669e-08 wk2=1.452943909e-07 pk2=-2.384048415e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.584068482e-01 ldsub=3.356002438e-11 wdsub=1.453258333e-10 pdsub=-2.185569740e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999992e-03 lcdscd=1.121188212e-18 wcdscd=5.664232972e-18 pcdscd=-8.422845754e-25 cit=0.0 voff='-2.075299990e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.569067098e-16 wvoff=-7.837899219e-16 pvoff=1.178749320e-22 nfactor=-6.134574575e+01 lnfactor=9.562494961e-06 wnfactor=4.141018107e-05 pnfactor=-6.227606441e-12 eta0=3.135593016e-02 leta0=-4.715649221e-09 weta0=-2.042029565e-08 peta0=3.071028683e-15 etab=-0.043998 u0=-3.036427888e-02 lu0=8.679390055e-09 wu0=3.434175851e-08 pu0=-5.244905546e-15 ua=4.331352307e-10 lua=-3.005085513e-16 wua=-7.517079844e-16 pua=1.551291363e-22 ub=-1.164158323e-17 lub=2.301733478e-24 wub=7.710124705e-24 pub=-1.332348938e-30 uc=1.576096325e-09 luc=-2.254499939e-16 wuc=-9.762718841e-16 puc=1.468225049e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.862244659e+06 lvsat=3.267682859e-01 wvsat=1.440624537e+00 pvsat=-2.251232183e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.690691819e-01 lketa=8.152232634e-08 wketa=3.530182181e-07 pketa=-5.309076284e-14 dwg=0.0 dwb=0.0 pclm=-1.047737130e+00 lpclm=1.540799100e-07 wpclm=8.904604567e-07 ppclm=-1.168246770e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.494484279e-07 lalpha0=5.706562851e-14 walpha0=2.471127531e-13 palpha0=-3.716353405e-20 alpha1=0.85 beta0=1.992691665e+01 lbeta0=-7.999607104e-07 wbeta0=-4.279469322e-06 pbeta0=5.805835024e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.686693084e-01 lkt1=3.010022753e-08 wkt1=1.710642403e-07 pkt1=-2.261255513e-14 kt2=-0.028878939 at=3.699275107e+05 lat=-4.755469050e-02 wat=-2.059272946e-01 pat=3.096961176e-8 ute=-2.397228847e+00 lute=1.906376330e-07 wute=6.216782825e-07 pute=-1.092473607e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.81 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.82 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.212001246e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.214741255e-06 wvth0=2.019659218e-08 pvth0=-4.039397405e-13 k1=7.466116614e-01 lk1=-3.572148663e-06 wk1=-7.528772312e-08 pk1=1.505783900e-12 k2=-1.130086766e-01 lk2=1.602877947e-06 wk2=3.717867333e-08 pk2=-7.435880035e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.343624387e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.217021741e-07 wvoff=1.835051541e-08 pvoff=-3.670174832e-13 nfactor=4.603746853e+00 lnfactor=-1.524323505e-05 wnfactor=-1.957574591e-07 pnfactor=3.915225724e-12 eta0=0.08 etab=-0.07 u0=8.025792333e-03 lu0=2.642473193e-07 wu0=6.011080706e-09 pu0=-1.202239644e-13 ua=-1.744751017e-09 lua=1.397228750e-14 wua=2.866357341e-16 pua=-5.732826756e-21 ub=1.493106929e-18 lub=-3.660410142e-24 wub=-7.516220008e-26 pub=1.503273390e-30 uc=6.585417669e-11 luc=-3.463503048e-16 wuc=-1.405229893e-18 puc=2.810514731e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.060004731e+00 la0=6.052023696e-06 wa0=1.857692258e-07 pa0=-3.715457153e-12 ags=5.476380673e-01 lags=-4.055240624e-06 wags=-1.273154529e-07 pags=2.546358838e-12 a1=0.0 a2=0.42385546 b0=1.112486784e-08 lb0=-2.221463796e-13 wb0=-7.225697527e-15 pb0=1.445167758e-19 b1=5.270682168e-08 lb1=-8.445929451e-13 wb1=-2.295181750e-14 pb1=4.590453242e-19 keta=-3.088153513e-02 lketa=5.267089995e-07 wketa=1.584211859e-08 pketa=-3.168485660e-13 dwg=0.0 dwb=0.0 pclm=-1.383881937e-01 lpclm=3.105324582e-06 wpclm=7.217304053e-08 ppclm=-1.443489030e-12 pdiblc1=0.39 pdiblc2=-7.048770547e-03 lpdiblc2=1.601850917e-07 wpdiblc2=4.264981571e-09 ppdiblc2=-8.530129902e-14 pdiblcb=1.055724067e+01 lpdiblcb=-2.116489510e-04 wpdiblcb=-5.939197917e-06 ppdiblcb=1.187862806e-10 drout=0.56 pscbe1=-4.923821975e+08 lpscbe1=1.434792445e+04 wpscbe1=2.342444857e+02 ppscbe1=-4.684981304e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.767420158e-01 lkt1=-1.927634528e-07 wkt1=-3.628146545e-09 pkt1=7.256434951e-14 kt2=-3.516743810e-02 lkt2=1.129923509e-07 wkt2=-1.768992198e-10 pkt2=3.538053564e-15 at=1.983344738e+05 lat=-4.666985988e-1 ute=-9.065670590e-01 lute=-4.176740474e-06 wute=-6.119112830e-08 pute=1.223846492e-12 ua1=5.688796016e-10 lua1=1.104262385e-14 wua1=2.585731307e-16 pua1=-5.171563715e-21 ub1=5.955929860e-20 lub1=-1.258083192e-23 wub1=-2.478782211e-25 pub1=4.957661342e-30 uc1=9.271776660e-11 luc1=-1.178011122e-15 wuc1=-1.307675531e-17 puc1=2.615402192e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.83 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.015346647e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.280055764e-07 wvth0=-5.438371812e-08 pvth0=1.927319028e-13 k1=5.828796647e-01 lk1=-2.262228669e-06 wk1=-8.212328385e-08 pk1=1.560471058e-12 k2=-4.330490943e-02 lk2=1.045220556e-06 wk2=3.520871719e-08 pk2=-7.278275841e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.095164997e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.229249466e-07 wvoff=-4.759647019e-09 pvoff=-1.821271477e-13 nfactor=1.112385167e+00 lnfactor=1.268902355e-05 wnfactor=1.461605283e-06 pnfactor=-9.344324244e-12 eta0=0.08 etab=-0.07 u0=5.568394788e-02 lu0=-1.170365595e-07 wu0=-1.821276292e-08 pu0=7.357625606e-14 ua=1.569307600e-09 lua=-1.254147723e-14 wua=-1.426035509e-15 pua=7.969212840e-21 ub=-1.048246406e-19 lub=9.123667207e-24 wub=8.511693887e-25 pub=-5.907741516e-30 uc=1.305103145e-10 luc=-8.636246876e-16 wuc=-6.791755487e-17 puc=5.602297534e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.120223562e+00 la0=-2.430141498e-06 wa0=-3.986023548e-07 pa0=9.597439822e-13 ags=2.586045904e-01 lags=-1.742859797e-06 wags=5.738331218e-08 pags=1.068696500e-12 a1=0.0 a2=0.42385546 b0=-7.638651043e-08 lb0=4.779788635e-13 wb0=4.974610383e-14 pb0=-3.112799110e-19 b1=-5.635028494e-08 lb1=2.790654916e-14 wb1=3.669767226e-14 pb1=-1.817391689e-20 keta=1.646582069e-02 lketa=1.479116402e-07 wketa=-1.907729573e-08 pketa=-3.747959796e-14 dwg=0.0 dwb=0.0 pclm=1.710465562e+00 lpclm=-1.168622836e-05 wpclm=-1.352374030e-06 ppclm=9.953444531e-12 pdiblc1=0.39 pdiblc2=3.176074161e-02 lpdiblc2=-1.503061801e-07 wpdiblc2=-1.875880237e-08 ppdiblc2=9.889797478e-14 pdiblcb=-3.177172200e+01 lpdiblcb=1.269993010e-04 wpdiblcb=1.781759375e-05 ppdiblcb=-7.127734168e-11 drout=0.56 pscbe1=1.644662413e+09 lpscbe1=-2.749268024e+03 wpscbe1=-5.645367612e+02 ppscbe1=1.705580995e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.224945882e-01 lkt1=1.732750160e-07 wkt1=2.034786643e-08 pkt1=-1.192531289e-13 kt2=-8.820774450e-02 lkt2=5.373355409e-07 wkt2=4.404533331e-08 pkt2=-3.502570976e-13 at=140000.0 ute=-3.105817286e+00 lute=1.341812125e-05 wute=1.052340334e-06 pute=-7.684840594e-12 ua1=-4.057530739e-10 lua1=1.884006633e-14 wua1=1.079396568e-15 pua1=-1.173847216e-20 ub1=-3.578449184e-19 lub1=-9.241434981e-24 wub1=-3.764207900e-25 pub1=5.986052153e-30 uc1=2.250531758e-10 luc1=-2.236746139e-15 wuc1=-1.664480834e-16 puc1=1.488570812e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.84 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='3.186852257e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.035027737e-07 wvth0=1.241739143e-07 pvth0=-5.215684430e-13 k1=-2.947195221e-01 lk1=1.248511219e-06 wk1=4.791800405e-07 pk1=-6.849617088e-13 k2=4.028066379e-01 lk2=-7.394000631e-07 wk2=-2.504518174e-07 pk2=4.149262475e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.311172409e+00 ldsub=7.485421266e-06 wdsub=1.218586062e-06 pdsub=-4.874820716e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.337536428e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.050289842e-06 wvoff=-2.083466135e-07 pvoff=6.323003205e-13 nfactor=1.204914533e+01 lnfactor=-3.106229338e-05 wnfactor=-5.551972836e-06 pnfactor=1.871273054e-11 eta0=-4.158606885e-01 leta0=1.983636635e-06 weta0=3.229253065e-07 peta0=-1.291827490e-12 etab=3.634882748e-01 letab=-1.734122593e-06 wetab=-2.823057711e-07 petab=1.129333466e-12 u0=3.445231451e-02 lu0=-3.210172439e-08 wu0=-3.800805021e-09 pu0=1.592278940e-14 ua=3.342584850e-09 lua=-1.963527959e-14 wua=-2.334296550e-15 pua=1.160261213e-20 ub=-5.136695914e-18 lub=2.925311976e-23 wub=3.794689634e-24 pub=-1.768297341e-29 uc=-2.454786209e-10 luc=6.404780657e-16 wuc=1.576871836e-16 puc=-3.422774119e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=8.527632932e-01 la0=2.640195154e-06 wa0=4.279537674e-07 pa0=-2.346803690e-12 ags=-1.038730269e+00 lags=3.446986900e-06 wags=7.658739492e-07 pags=-1.765543068e-12 a1=0.0 a2=0.42385546 b0=2.121750412e-07 lb0=-6.763801704e-13 wb0=-1.381772982e-13 pb0=4.404871750e-19 b1=3.634657342e-08 lb1=-3.429171288e-13 wb1=-2.367041517e-14 pb1=2.233220368e-19 keta=2.022048610e-01 lketa=-5.951171451e-07 wketa=-1.132105954e-07 pketa=3.390904068e-13 dwg=0.0 dwb=0.0 pclm=-3.299953641e+00 lpclm=8.357407523e-06 wpclm=2.480697326e-06 ppclm=-5.380339624e-12 pdiblc1=0.39 pdiblc2=-5.177636595e-03 lpdiblc2=-2.538224350e-09 wpdiblc2=4.278413787e-09 ppdiblc2=6.740102616e-15 pdiblcb=5.296551706e-02 lpdiblcb=-3.118925527e-07 wpdiblcb=-5.077441926e-08 ppdiblcb=2.031175298e-13 drout=0.56 pscbe1=1.114855946e+09 lpscbe1=-6.298350007e+02 wpscbe1=-2.763933918e+02 ppscbe1=5.528948534e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-5.295150438e-01 lkt1=1.001437783e-06 wkt1=1.522438686e-07 pkt1=-6.468887090e-13 kt2=-8.070923640e-02 lkt2=5.073385766e-07 wkt2=3.712774665e-08 pkt2=-3.225840461e-13 at=1.573914787e+05 lat=-6.957271488e-02 wat=7.433374980e-03 pat=-2.973640637e-8 ute=-7.238503639e+00 lute=2.995048254e-05 wute=3.575216997e-06 pute=-1.777733369e-11 ua1=-1.850064234e-08 lua1=9.122669848e-14 wua1=1.159244689e-14 pua1=-5.379478406e-20 ub1=1.540798430e-17 lub1=-7.231091630e-23 wub1=-9.487277020e-24 pub1=4.243303942e-29 uc1=-9.659102569e-11 luc1=-9.500435698e-16 wuc1=5.877014636e-17 puc1=5.876098329e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.85 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='8.042249147e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.776645031e-08 wvth0=-1.776040530e-07 pvth0=8.210548677e-14 k1=6.468961762e-01 lk1=-6.350883493e-07 wk1=-3.080091740e-08 pk1=3.351996097e-13 k2=-8.862583514e-02 lk2=2.436570332e-07 wk2=2.450273140e-08 pk2=-1.350903573e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.602462119e+00 ldsub=-4.344160021e-06 wdsub=-2.437172124e-06 pdsub=2.438125059e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.272737657e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.198433681e-08 wvoff=1.477845971e-07 pvoff=-8.010134797e-14 nfactor=-4.931803891e+00 lnfactor=2.906244616e-06 wnfactor=5.038704115e-06 pnfactor=-2.472764314e-12 eta0=1.149220055e+00 leta0=-1.147136799e-06 weta0=-6.458504098e-07 peta0=6.461027342e-13 etab=-9.225959290e-01 letab=8.385486734e-07 wetab=5.646115422e-07 petab=-5.648323053e-13 u0=9.801978587e-03 lu0=1.720858573e-08 wu0=1.138950525e-08 pu0=-1.446377056e-14 ua=-9.929291739e-09 lua=6.913662895e-15 wua=5.868036349e-15 pua=-4.805260774e-21 ub=1.412986726e-17 lub=-9.287539806e-24 wub=-8.192934820e-24 pub=6.296962656e-30 uc=-1.115873300e-10 luc=3.726431323e-16 wuc=9.744211970e-17 puc=-2.217637283e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.892206602e+04 lvsat=1.021758394e-01 wvsat=2.674912952e-02 pvsat=-5.350871796e-8 a0=6.999550514e+00 la0=-9.655782680e-06 wa0=-3.653735593e-06 pa0=5.818170971e-12 ags=4.314892342e+00 lags=-7.262351590e-06 wags=-2.588613558e-06 pags=4.944743552e-12 a1=0.0 a2=0.42385546 b0=2.500992201e-07 lb0=-7.522433566e-13 wb0=-1.628751163e-13 pb0=4.898924681e-19 b1=-2.001955281e-07 lb1=1.302595623e-13 wb1=1.303757361e-13 pb1=-8.483049788e-20 keta=-6.506983864e-01 lketa=1.111022835e-06 wketa=4.060268569e-07 pketa=-6.995875195e-13 dwg=0.0 dwb=0.0 pclm=2.203217795e+00 lpclm=-2.651087090e-06 wpclm=-1.157516946e-06 ppclm=1.897511462e-12 pdiblc1=5.390330599e-01 lpdiblc1=-2.981243917e-07 wpdiblc1=-6.363782049e-08 ppdiblc1=1.273005234e-13 pdiblc2=-2.564189589e-02 lpdiblc2=3.839829577e-08 wpdiblc2=1.981654525e-08 ppdiblc2=-2.434223571e-14 pdiblcb=1.502650000e-01 lpdiblcb=-5.065295627e-07 wpdiblcb=-9.826130131e-08 ppdiblcb=2.981098613e-13 drout=3.981758719e+00 ldrout=-6.844855346e-06 wdrout=-2.122394365e-06 pdrout=4.245618587e-12 pscbe1=3.876199809e+08 lpscbe1=8.249212788e+02 wpscbe1=2.685591884e+02 ppscbe1=-5.372233835e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.428783480e-05 lalpha0=-6.852906442e-11 walpha0=-2.230935906e-11 palpha0=4.462744108e-17 alpha1=1.957544281e+00 lalpha1=-2.215521611e-06 walpha1=-6.216003671e-07 palpha1=1.243443780e-12 beta0=3.634341167e+01 lbeta0=-4.497561435e-05 wbeta0=-1.464214198e-05 pbeta0=2.929000904e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=8.654253384e-02 lkt1=-2.309182505e-07 wkt1=-2.691428415e-07 pkt1=1.960494734e-13 kt2=4.389055626e-01 lkt2=-5.320941908e-07 wkt2=-2.852889709e-07 pkt2=3.223754538e-13 at=1.587042509e+04 lat=2.135247271e-01 wat=7.868601478e-02 pat=-1.722695458e-7 ute=1.634436459e+01 lute=-1.722447482e-05 wute=-1.051251800e-05 pute=1.040364461e-11 ua1=5.319138333e-08 lua1=-5.218538443e-14 wua1=-3.074862473e-14 pua1=3.090391454e-20 ub1=-4.011353472e-17 lub1=3.875383065e-23 wub1=2.305923212e-23 pub1=-2.267270454e-29 uc1=-1.018027742e-09 luc1=8.931901437e-16 wuc1=6.118569544e-16 puc1=-5.187800402e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.86 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='8.857756556e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.493490775e-07 wvth0=-1.911360188e-07 pvth0=9.564274357e-14 k1=-4.512339609e-01 lk1=4.634711567e-07 wk1=6.087732982e-07 pk1=-3.046246795e-13 k2=3.192061816e-01 lk2=-1.643344459e-07 wk2=-2.211560907e-07 pk2=1.106645174e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615564e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.670860321e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.118121698e-07 wvoff=1.354820659e-07 pvoff=-6.779400644e-14 nfactor=-7.102416557e+00 lnfactor=5.077705992e-06 wnfactor=5.135819868e-06 pnfactor=-2.569918039e-12 eta0=-4.853179767e-01 leta0=4.880403377e-07 weta0=-4.062747498e-13 peta0=2.032962284e-19 etab=-1.681904925e-01 letab=8.384826436e-8 u0=3.454176684e-02 lu0=-7.540875777e-09 wu0=-6.139624018e-09 pu0=3.072212602e-15 ua=-4.593839643e-09 lua=1.576124638e-15 wua=2.130139953e-15 pua=-1.065902861e-21 ub=8.111606463e-18 lub=-3.266925871e-24 wub=-3.798351203e-24 pub=1.900660757e-30 uc=4.694462594e-10 luc=-2.086176412e-16 wuc=-2.485670174e-16 puc=1.243806984e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-2.394417634e+04 lvsat=1.550627525e-01 wvsat=-5.349825905e-02 pvsat=2.677004734e-8 a0=-6.692673442e+00 la0=4.041794935e-06 wa0=4.326013535e-06 pa0=-2.164698239e-12 ags=-6.047916438e+00 lags=3.104509048e-06 wags=4.710235692e-06 pags=-2.356959548e-12 a1=0.0 a2=0.42385546 b0=-1.004092695e-06 lb0=5.024389480e-13 wb0=6.539073352e-13 pb0=-3.272093454e-19 b1=-1.400284845e-07 lb1=7.006899341e-14 wb1=9.119243033e-14 pb1=-4.563187140e-20 keta=9.272589265e-01 lketa=-4.675514593e-07 wketa=-5.868038123e-07 pketa=2.936313465e-13 dwg=0.0 dwb=0.0 pclm=-1.346178989e+00 lpclm=8.996975080e-07 wpclm=1.479083854e-06 ppclm=-7.401202487e-13 pdiblc1=4.491812363e-01 lpdiblc1=-2.082374361e-07 wpdiblc1=1.272756410e-07 ppdiblc1=-6.368758526e-14 pdiblc2=2.544627381e-02 lpdiblc2=-1.270984941e-08 wpdiblc2=-9.035884392e-09 ppdiblc2=4.521475227e-15 pdiblcb=-6.177324269e-01 lpdiblcb=2.617681512e-07 wpdiblcb=3.996202797e-07 ppdiblcb=-1.999663914e-13 drout=-6.723861418e+00 ldrout=3.864950689e-06 wdrout=4.244788731e-06 pdrout=-2.124054078e-12 pscbe1=1.988096935e+09 lpscbe1=-7.761814621e+02 wpscbe1=-5.371183768e+02 ppscbe1=2.687692017e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-7.235869595e-05 lalpha0=3.815916513e-11 walpha0=4.461871812e-11 palpha0=-2.232680498e-17 alpha1=-1.365088561e+00 lalpha1=1.108410380e-06 walpha1=1.243200734e-06 palpha1=-6.220864586e-13 beta0=-3.526807489e+01 lbeta0=2.666387230e-05 wbeta0=2.928428396e-05 pbeta0=-1.465359214e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-9.516038467e-03 lkt1=-1.348221193e-07 wkt1=-1.463972058e-07 pkt1=7.325584422e-14 kt2=-1.492867183e-01 lkt2=5.632807329e-08 wkt2=7.394986993e-08 pkt2=-3.700384937e-14 at=4.481391226e+05 lat=-2.189129874e-01 wat=-1.871055295e-01 pat=9.362592300e-8 ute=-4.361356291e-01 lute=-4.374134255e-07 wute=-2.259675782e-07 pute=1.130721424e-13 ua1=1.221273519e-09 lua1=-1.949543095e-16 wua1=2.865342053e-16 pua1=-1.433791375e-22 ub1=-2.118403788e-18 lub1=7.438436252e-25 wub1=7.910874670e-25 pub1=-3.958530487e-31 uc1=-2.562162105e-10 luc1=1.310807443e-16 wuc1=1.866323007e-16 puc1=-9.338912356e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.87 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.303289752e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.152585767e-8 k1=4.221882219e-02 lk1=2.165518251e-7 k2=1.272986658e-01 lk2=-6.830565219e-08 wk2=-2.775557562e-23 pk2=6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383648e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267778e-8 nfactor=4.152229107e+00 lnfactor=-5.540174069e-7 eta0=9.800711344e-01 leta0=-2.452271850e-7 etab=4.281583539e-02 letab=-2.173740306e-08 wetab=1.387778781e-23 petab=-5.421010862e-30 u0=1.871952528e-02 lu0=3.764314976e-10 ua=-1.777587834e-09 lua=1.668975788e-16 ub=1.993952344e-18 lub=-2.057068089e-25 wub=-1.540743956e-39 uc=1.245140400e-11 luc=2.005847147e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.384900615e+05 lvsat=-2.629607820e-2 a0=1.269019515e+00 la0=5.783543445e-8 ags=-9.392106230e-01 lags=5.481586371e-07 wags=-2.220446049e-22 pags=1.110223025e-28 a1=0.0 a2=0.42385546 b0=-4.603925132e-17 lb0=1.152781418e-23 b1=1.027396975e-17 lb1=-2.572509561e-24 keta=6.904029211e-02 lketa=-3.810657865e-08 wketa=2.081668171e-23 pketa=-1.040834086e-29 dwg=0.0 dwb=0.0 pclm=6.653835068e-01 lpclm=-1.068702608e-07 wpclm=-4.440892099e-22 pdiblc1=-2.914152067e-01 lpdiblc1=1.623503586e-07 ppdiblc1=-1.387778781e-29 pdiblc2=-8.326311299e-03 lpdiblc2=4.189648227e-09 wpdiblc2=3.089976192e-24 ppdiblc2=1.151964808e-30 pdiblcb=-8.590105794e-02 lpdiblcb=-4.355479349e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974521e+07 lpscbe1=1.776524482e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465818e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-8 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438220939e+03 lat=9.053815040e-3 ute=-1.301500893e+00 lute=-4.392435834e-9 ua1=1.688524505e-09 lua1=-4.287624978e-16 ub1=-1.973606354e-18 lub1=6.713882924e-25 wub1=7.703719778e-40 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=4.523643975e-32 puc1=3.231174268e-39 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.88 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.724931888e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322408849e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232527937e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767236523e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665325738e-16 ags=1.250000000e+00 lags=5.706635164e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.562972222e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223438018e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387523651e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448147158e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435282e-25 ub1=7.077531678e-19 lub1=3.881557729e-34 uc1=1.471862500e-10 luc1=-5.620278672e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.89 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='8.324779087e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.020461593e-08 wvth0=-1.078769616e-07 pvth0=1.946003298e-14 k1=0.90707349 k2=-9.227639866e-02 lk2=-8.991402185e-09 wk2=-1.671609289e-08 pk2=3.015432712e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999998e-03 lcdscd=4.032121859e-19 wcdscd=2.077199523e-18 pcdscd=-3.747080771e-25 cit=0.0 voff='-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.409361599e-17 nfactor=2.246464102e+00 lnfactor=-1.201078162e-09 wnfactor=-3.736857242e-09 pnfactor=6.740954148e-16 eta0=1.493096587e-09 leta0=-2.245188128e-16 weta0=5.416137448e-19 peta0=-9.770224504e-26 etab=-0.043998 u0=-8.472696194e-02 lu0=1.994473923e-08 wu0=6.974502095e-08 pu0=-1.258137407e-14 ua=1.432666132e-09 lua=-4.508294850e-16 wua=-1.402644488e-15 pua=2.530244418e-22 ub=-8.647940787e-18 lub=1.851517514e-24 wub=5.760539011e-24 pub=-1.039149393e-30 uc=7.700399984e-11 luc=2.365891648e-26 wuc=-1.422750654e-28 puc=2.569429778e-35 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.113256855e+06 lvsat=-1.566220151e-01 wvsat=-4.971470199e-01 pvsat=8.968084806e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000008e-02 lketa=1.270780703e-17 wketa=8.137934771e-20 pketa=-1.468269950e-26 dwg=0.0 dwb=0.0 pclm=1.194459649e+00 lpclm=-1.831263154e-07 wpclm=-5.697522582e-07 ppclm=1.027781796e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.832266417e-24 walpha0=-1.628420841e-25 palpha0=2.938145536e-32 alpha1=0.85 beta0=1.019114168e+01 lbeta0=6.623943411e-07 wbeta0=2.060876241e-06 pbeta0=-3.717635260e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.621629336e-02 lkt1=-3.344469693e-08 wkt1=-1.040549061e-07 pkt1=1.877056856e-14 kt2=-0.028878939 at=5.372048691e+04 lat=1.395307481e-11 wat=-3.469176590e-14 pat=6.257323548e-21 ute=-2.233757785e+00 lute=1.655985860e-07 wute=5.152190612e-07 pute=-9.294088166e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.90 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.91 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-6 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-7 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 pb0=-9.926167351e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-07 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-08 wkt1=-1.776356839e-21 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344737e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 wuc1=-2.067951531e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.92 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-07 pk2=4.440892099e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008797e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539118e-02 lketa=8.113189461e-8 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=-1.776356839e-21 ppclm=7.105427358e-27 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-08 ppdiblc2=-5.551115123e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 uc1=-7.151779256e-11 luc1=4.155336487e-16 wuc1=-2.067951531e-31 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.93 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155423e-01 leta0=-3.180932596e-7 etab=-1.395135872e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 wb0=5.293955920e-29 b1=-5.828486835e-09 lb1=5.498972206e-14 keta=4.904572511e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-6 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-08 wpdiblcb=-2.220446049e-22 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-1 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 ub1=-1.496090981e-18 lub1=3.294685946e-24 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.94 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-09 peta0=1.040834086e-29 etab=8.340779512e-02 letab=-1.678483982e-07 wetab=-2.220446049e-22 petab=-4.267419751e-28 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 pua=-3.308722450e-36 ub=-4.679975144e-19 lub=1.932152691e-24 uc=6.203139367e-11 luc=-2.248718272e-17 wuc=-4.135903063e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024581e-01 lags=1.548007492e-06 pags=-3.552713679e-27 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 pb0=2.117582368e-34 b1=3.210308126e-08 lb1=-2.088824537e-14 keta=7.274507804e-02 lketa=-1.354760365e-07 wketa=1.110223025e-22 pketa=3.885780586e-28 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-09 wpdiblc2=5.551115123e-23 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=-4.235164736e-27 palpha0=1.482307658e-32 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-08 wkt2=-4.440892099e-22 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-06 wute=-1.421085472e-20 ua1=-1.595365930e-09 lua1=2.878054409e-15 pua1=3.308722450e-36 ub1=9.725424449e-19 lub1=-1.643546140e-24 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.95 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.452166476e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.106358502e-8 k1=6.334555282e-01 lk1=-7.929770144e-8 k2=-7.484146749e-02 lk2=3.284345126e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615564e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891553e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980654741e-9 nfactor=2.048395157e+00 lnfactor=4.987221675e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-4.440892099e-22 peta0=-5.828670879e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.360241444e-02 lu0=-2.066922291e-9 ua=-7.984359621e-10 lua=-3.230612055e-16 ub=1.343846382e-18 lub=1.196003632e-25 uc=2.655884652e-11 luc=1.299923420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.192653730e+05 lvsat=2.027606214e-01 pvsat=4.656612873e-22 a0=1.015255643e+00 la0=1.848165925e-7 ags=2.344605312e+00 lags=-1.095033302e-6 a1=0.0 a2=0.42385546 b0=1.610149323e-07 lb0=-8.057042298e-14 b1=2.245477638e-08 lb1=-1.123616801e-14 keta=-1.182861545e-01 lketa=5.562988931e-8 dwg=0.0 dwb=0.0 pclm=1.289197291e+00 lpclm=-4.190210639e-7 pdiblc1=6.759562121e-01 lpdiblc1=-3.217135930e-7 pdiblc2=9.346473028e-03 lpdiblc2=-4.653653995e-9 pdiblcb=9.429603789e-02 lpdiblcb=-9.452448433e-08 wpdiblcb=1.734723476e-22 ppdiblcb=-2.029626467e-28 drout=8.393443483e-01 ldrout=8.039059217e-8 pscbe1=1.031079505e+09 lpscbe1=-2.972985529e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266840e-06 lalpha0=-1.621900755e-12 alpha1=0.85 beta0=1.690956677e+01 lbeta0=5.546500095e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611032e-01 lkt1=-4.297596482e-9 kt2=-1.752560647e-02 lkt2=-9.604001224e-9 at=1.147614896e+05 lat=-5.209382031e-2 ute=-8.387562066e-01 lute=-2.359457121e-7 ua1=1.731809447e-09 lua1=-4.504218931e-16 ub1=-7.088737332e-19 lub1=3.852747156e-26 uc1=7.631824104e-11 luc1=-3.531650240e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.96 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.303289752e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.152585767e-8 k1=4.221882219e-02 lk1=2.165518251e-7 k2=1.272986658e-01 lk2=-6.830565219e-08 wk2=-1.110223025e-22 pk2=1.942890293e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383648e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267778e-8 nfactor=4.152229107e+00 lnfactor=-5.540174069e-7 eta0=9.800711344e-01 leta0=-2.452271850e-7 etab=4.281583539e-02 letab=-2.173740306e-08 wetab=-4.857225733e-23 petab=4.683753385e-29 u0=1.871952528e-02 lu0=3.764314976e-10 ua=-1.777587834e-09 lua=1.668975788e-16 ub=1.993952344e-18 lub=-2.057068089e-25 uc=1.245140400e-11 luc=2.005847147e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.384900615e+05 lvsat=-2.629607820e-2 a0=1.269019515e+00 la0=5.783543445e-8 ags=-9.392106230e-01 lags=5.481586371e-07 wags=1.776356839e-21 pags=-1.776356839e-27 a1=0.0 a2=0.42385546 b0=-4.603925132e-17 lb0=1.152781418e-23 b1=1.027396975e-17 lb1=-2.572509561e-24 keta=6.904029211e-02 lketa=-3.810657865e-08 wketa=-1.110223025e-22 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=6.653835068e-01 lpclm=-1.068702608e-7 pdiblc1=-2.914152067e-01 lpdiblc1=1.623503586e-07 wpdiblc1=-4.440892099e-22 ppdiblc1=3.330669074e-28 pdiblc2=-8.326311299e-03 lpdiblc2=4.189648227e-09 wpdiblc2=2.125036258e-23 ppdiblc2=6.179952383e-30 pdiblcb=-8.590105794e-02 lpdiblcb=-4.355479349e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974521e+07 lpscbe1=1.776524482e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465818e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-8 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438220939e+03 lat=9.053815040e-03 pat=-2.910383046e-23 ute=-1.301500893e+00 lute=-4.392435834e-9 ua1=1.688524505e-09 lua1=-4.287624978e-16 ub1=-1.973606354e-18 lub1=6.713882924e-25 pub1=-1.540743956e-45 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=-1.033975766e-31 puc1=1.550963649e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.97 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.725464795e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322320031e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232475895e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.766986723e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665316856e-16 ags=1.250000000e+00 lags=5.706368711e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.563105449e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223465773e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387237549e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448174913e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732436057e-25 ub1=7.077531678e-19 lub1=3.881534617e-34 uc1=1.471862500e-10 luc1=-5.619865082e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.98 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='-5.678691211e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.024053851e-07 wvth0=6.780566061e-07 pvth0=-1.223153092e-13 k1=0.90707349 k2=-1.367273487e+00 lk2=2.210065975e-07 wk2=6.988658227e-07 pk2=-1.260691046e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000026e-03 lcdscd=-4.702474521e-18 wcdscd=-1.380795478e-17 pcdscd=2.490826989e-24 cit=0.0 voff='-2.075300002e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.409272781e-17 nfactor=2.246463368e+00 lnfactor=-1.200945814e-09 wnfactor=-3.736445473e-09 pnfactor=6.740211354e-16 eta0=1.493096730e-09 leta0=-2.245188117e-16 weta0=5.416171744e-19 peta0=-9.770286371e-26 etab=-0.043998 u0=9.451685443e-01 lu0=-1.658391410e-07 wu0=-5.082755928e-07 pu0=9.168834245e-14 ua=1.432519508e-09 lua=-4.508030353e-16 wua=-1.402562196e-15 pua=2.530095971e-22 ub=-8.647861908e-18 lub=1.851503285e-24 wub=5.760494741e-24 pub=-1.039141407e-30 uc=7.700399984e-11 luc=2.400891728e-26 wuc=9.462946208e-28 puc=-1.708127965e-34 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.085396075e+07 lvsat=2.002156336e+00 wvsat=6.219358124e+00 pvsat=-1.121916231e-6 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000008e-02 lketa=1.250688442e-17 wketa=-5.426770144e-19 pketa=9.803269307e-26 dwg=0.0 dwb=0.0 pclm=1.194459627e+00 lpclm=-1.831263114e-07 wpclm=-5.697522456e-07 ppclm=1.027781773e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.430984559e-24 walpha0=1.085896238e-24 palpha0=-1.958763691e-31 alpha1=0.85 beta0=1.023373151e+01 lbeta0=6.547115191e-07 wbeta0=2.036973040e-06 pbeta0=-3.674516037e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-5.014731662e-02 lkt1=-3.273557571e-08 wkt1=-1.018486507e-07 pkt1=1.837257995e-14 kt2=-0.028878939 at=5.372048691e+04 lat=1.403875649e-11 wat=2.328306437e-13 pat=-4.190951586e-20 ute=-2.223110315e+00 lute=1.636778782e-07 wute=5.092432536e-07 pute=-9.186289976e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.99 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.100 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-6 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-7 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 wb0=-5.169878828e-31 pb0=2.192028623e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-7 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+03 ppscbe1=-3.814697266e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-8 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344738e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.101 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-07 pk2=1.110223025e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008797e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 wb0=-6.617444900e-30 pb0=-2.646977960e-35 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539118e-02 lketa=8.113189461e-8 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=4.440892099e-22 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-08 ppdiblc2=-1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 uc1=-7.151779256e-11 luc1=4.155336487e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.102 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155423e-01 leta0=-3.180932596e-7 etab=-1.395135872e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 wb0=-2.646977960e-29 pb0=-1.058791184e-34 b1=-5.828486835e-09 lb1=5.498972206e-14 keta=4.904572511e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-06 wpclm=1.776356839e-21 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-8 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-1 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 ub1=-1.496090981e-18 lub1=3.294685946e-24 pub1=-3.081487911e-45 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.103 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-9 etab=8.340779513e-02 letab=-1.678483982e-07 wetab=-5.204170428e-23 petab=6.938893904e-29 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 ub=-4.679975144e-19 lub=1.932152691e-24 pub=-1.540743956e-45 uc=6.203139367e-11 luc=-2.248718272e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024581e-01 lags=1.548007492e-6 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 pb0=5.293955920e-35 b1=3.210308126e-08 lb1=-2.088824537e-14 wb1=5.293955920e-29 keta=7.274507804e-02 lketa=-1.354760365e-07 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-9 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=1.058791184e-28 palpha0=-1.164670302e-33 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-08 wkt2=1.110223025e-22 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-6 ua1=-1.595365930e-09 lua1=2.878054409e-15 wua1=1.240770919e-30 pua1=8.271806126e-37 ub1=9.725424449e-19 lub1=-1.643546140e-24 wub1=3.851859889e-40 pub1=-1.155557967e-45 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.104 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.452166476e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.106358502e-8 k1=6.334555282e-01 lk1=-7.929770144e-8 k2=-7.484146749e-02 lk2=3.284345126e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615564e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891553e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980654741e-9 nfactor=2.048395157e+00 lnfactor=4.987221675e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-3.191891196e-22 peta0=-2.255140519e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.360241444e-02 lu0=-2.066922291e-9 ua=-7.984359621e-10 lua=-3.230612055e-16 ub=1.343846382e-18 lub=1.196003632e-25 uc=2.655884652e-11 luc=1.299923420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.192653730e+05 lvsat=2.027606214e-1 a0=1.015255643e+00 la0=1.848165925e-7 ags=2.344605312e+00 lags=-1.095033302e-6 a1=0.0 a2=0.42385546 b0=1.610149323e-07 lb0=-8.057042298e-14 b1=2.245477638e-08 lb1=-1.123616801e-14 keta=-1.182861545e-01 lketa=5.562988931e-8 dwg=0.0 dwb=0.0 pclm=1.289197291e+00 lpclm=-4.190210639e-7 pdiblc1=6.759562121e-01 lpdiblc1=-3.217135930e-07 ppdiblc1=-4.440892099e-28 pdiblc2=9.346473028e-03 lpdiblc2=-4.653653995e-9 pdiblcb=9.429603789e-02 lpdiblcb=-9.452448433e-08 wpdiblcb=4.900593820e-23 ppdiblcb=4.987329993e-29 drout=8.393443483e-01 ldrout=8.039059217e-8 pscbe1=1.031079505e+09 lpscbe1=-2.972985529e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266840e-06 lalpha0=-1.621900755e-12 alpha1=0.85 beta0=1.690956677e+01 lbeta0=5.546500095e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611032e-01 lkt1=-4.297596482e-9 kt2=-1.752560647e-02 lkt2=-9.604001224e-9 at=1.147614896e+05 lat=-5.209382031e-2 ute=-8.387562066e-01 lute=-2.359457121e-7 ua1=1.731809447e-09 lua1=-4.504218931e-16 ub1=-7.088737332e-19 lub1=3.852747156e-26 uc1=7.631824104e-11 luc1=-3.531650240e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.105 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.303289752e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.152585767e-8 k1=4.221882219e-02 lk1=2.165518251e-7 k2=1.272986658e-01 lk2=-6.830565219e-08 wk2=-5.551115123e-23 pk2=-4.163336342e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383648e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267778e-8 nfactor=4.152229107e+00 lnfactor=-5.540174069e-07 wnfactor=-7.105427358e-21 eta0=9.800711344e-01 leta0=-2.452271850e-7 etab=4.281583539e-02 letab=-2.173740306e-08 wetab=1.387778781e-23 petab=8.673617380e-30 u0=1.871952528e-02 lu0=3.764314976e-10 ua=-1.777587834e-09 lua=1.668975788e-16 ub=1.993952344e-18 lub=-2.057068089e-25 uc=1.245140400e-11 luc=2.005847147e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.384900615e+05 lvsat=-2.629607820e-2 a0=1.269019515e+00 la0=5.783543445e-8 ags=-9.392106230e-01 lags=5.481586371e-07 wags=-4.440892099e-22 pags=-1.110223025e-28 a1=0.0 a2=0.42385546 b0=-4.603925132e-17 lb0=1.152781418e-23 b1=1.027396975e-17 lb1=-2.572509561e-24 keta=6.904029211e-02 lketa=-3.810657865e-08 wketa=-5.551115123e-23 pketa=6.938893904e-30 dwg=0.0 dwb=0.0 pclm=6.653835068e-01 lpclm=-1.068702608e-7 pdiblc1=-2.914152067e-01 lpdiblc1=1.623503586e-07 wpdiblc1=-1.110223025e-22 ppdiblc1=5.551115123e-29 pdiblc2=-8.326311299e-03 lpdiblc2=4.189648227e-09 wpdiblc2=-2.168404345e-25 ppdiblc2=-2.602085214e-30 pdiblcb=-8.590105794e-02 lpdiblcb=-4.355479349e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974521e+07 lpscbe1=1.776524482e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465818e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-8 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438220939e+03 lat=9.053815040e-03 pat=7.275957614e-24 ute=-1.301500893e+00 lute=-4.392435834e-9 ua1=1.688524505e-09 lua1=-4.287624978e-16 ub1=-1.973606354e-18 lub1=6.713882924e-25 wub1=-1.540743956e-39 pub1=-3.851859889e-46 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=-3.877409121e-32 puc1=9.693522803e-39 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.106 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.725109524e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322408849e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232545284e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767208767e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665316856e-16 ags=1.250000000e+00 lags=5.706723982e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.562927813e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223451895e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416724598e-16 pscbe1=7.914198799e+08 lpscbe1=2.387619019e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448174913e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435540e-25 ub1=7.077531678e-19 lub1=3.881534617e-34 uc1=1.471862500e-10 luc1=-5.620278672e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.107 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.056294159e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.679501053e-08 wvth0=1.414233256e-07 pvth0=-2.551149513e-14 k1=0.90707349 k2=2.096955826e-01 lk2=-6.346442986e-08 wk2=-1.704257609e-07 pk2=3.074327344e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585017754e-01 ldsub=2.313056177e-11 wdsub=7.068277868e-11 pdsub=-1.275053713e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.839153829e-19 cit=0.0 voff='-5.767404296e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.660223861e-08 wvoff=2.035242956e-07 pvoff=-3.671395120e-14 nfactor=-1.428319278e+01 lnfactor=2.980600256e-06 wnfactor=9.108104269e-06 pnfactor=-1.643020037e-12 eta0=1.783339662e-02 leta0=-3.216983883e-09 weta0=-9.830515412e-09 peta0=1.773336506e-15 etab=-0.043998 u0=-2.986511643e-01 lu0=5.853474002e-08 wu0=1.773700710e-07 pu0=-3.199596449e-14 ua=-6.409135178e-10 lua=-7.677437833e-17 wua=-2.595988281e-16 pua=4.682929220e-23 ub=2.506645255e-17 lub=-4.230255614e-24 wub=-1.282425139e-23 pub=2.313379532e-30 uc=3.495542053e-10 luc=-4.916560408e-17 wuc=-1.502411203e-16 puc=2.710214594e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.606406842e+06 lvsat=-1.508318834e+00 wvsat=-4.508013829e+00 pvsat=8.132051226e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000008e-02 lketa=1.268474215e-17 dwg=0.0 dwb=0.0 pclm=-3.426700006e-01 lpclm=9.415803923e-08 wpclm=2.775781644e-07 ppclm=-5.007260265e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.786314880e-24 alpha1=0.85 beta0=1.392897432e+01 lbeta0=-1.187702761e-8 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.918229625e-01 lkt1=4.693873573e-08 wkt1=1.416215157e-07 pkt1=-2.554724684e-14 kt2=-0.028878939 at=5.372048691e+04 lat=1.396285370e-11 ute=3.619587319e-01 lute=-3.026453122e-07 wute=-9.157553778e-07 pute=1.651940284e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.108 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.109 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-6 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-07 wags=-1.776356839e-21 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 wb0=1.137373342e-30 pb0=-5.128519798e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-7 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-8 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344738e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.110 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-07 pk2=-4.440892099e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008797e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 pb0=-1.058791184e-34 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539118e-02 lketa=8.113189461e-08 wketa=-5.551115123e-23 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=-1.776356839e-21 ppclm=5.329070518e-27 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-08 ppdiblc2=5.551115123e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 uc1=-7.151779256e-11 luc1=4.155336487e-16 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.111 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155422e-01 leta0=-3.180932596e-7 etab=-1.395135873e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 wb0=5.293955920e-29 pb0=1.058791184e-34 b1=-5.828486835e-09 lb1=5.498972206e-14 pb1=-1.058791184e-34 keta=4.904572512e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-6 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-8 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-1 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 ub1=-1.496090981e-18 lub1=3.294685946e-24 pub1=-1.232595164e-44 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.112 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-09 peta0=-3.469446952e-30 etab=8.340779513e-02 letab=-1.678483982e-07 wetab=-2.012279232e-22 petab=3.365363543e-28 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 pua=3.308722450e-36 ub=-4.679975144e-19 lub=1.932152691e-24 pub=-3.081487911e-45 uc=6.203139367e-11 luc=-2.248718272e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024581e-01 lags=1.548007492e-06 pags=-3.552713679e-27 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 b1=3.210308126e-08 lb1=-2.088824537e-14 keta=7.274507804e-02 lketa=-1.354760365e-07 wketa=-1.110223025e-22 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-09 wpdiblc2=-5.551115123e-23 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=-1.270549421e-27 palpha0=1.905824131e-33 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-8 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-6 ua1=-1.595365930e-09 lua1=2.878054409e-15 pua1=-1.654361225e-36 ub1=9.725424449e-19 lub1=-1.643546140e-24 wub1=-1.540743956e-39 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.113 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.452166476e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.106358502e-8 k1=6.334555282e-01 lk1=-7.929770144e-8 k2=-7.484146749e-02 lk2=3.284345126e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615564e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891553e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980654741e-9 nfactor=2.048395157e+00 lnfactor=4.987221675e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=6.938893904e-22 peta0=6.245004514e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.360241444e-02 lu0=-2.066922291e-9 ua=-7.984359621e-10 lua=-3.230612055e-16 ub=1.343846382e-18 lub=1.196003632e-25 uc=2.655884652e-11 luc=1.299923420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.192653730e+05 lvsat=2.027606214e-01 pvsat=4.656612873e-22 a0=1.015255643e+00 la0=1.848165925e-7 ags=2.344605312e+00 lags=-1.095033302e-6 a1=0.0 a2=0.42385546 b0=1.610149323e-07 lb0=-8.057042298e-14 b1=2.245477638e-08 lb1=-1.123616801e-14 keta=-1.182861545e-01 lketa=5.562988931e-8 dwg=0.0 dwb=0.0 pclm=1.289197291e+00 lpclm=-4.190210639e-7 pdiblc1=6.759562121e-01 lpdiblc1=-3.217135930e-7 pdiblc2=9.346473028e-03 lpdiblc2=-4.653653995e-9 pdiblcb=9.429603789e-02 lpdiblcb=-9.452448433e-08 wpdiblcb=-4.163336342e-23 ppdiblcb=-1.873501354e-28 drout=8.393443483e-01 ldrout=8.039059217e-8 pscbe1=1.031079505e+09 lpscbe1=-2.972985529e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266840e-06 lalpha0=-1.621900755e-12 alpha1=0.85 beta0=1.690956677e+01 lbeta0=5.546500095e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611032e-01 lkt1=-4.297596482e-9 kt2=-1.752560647e-02 lkt2=-9.604001224e-9 at=1.147614896e+05 lat=-5.209382031e-2 ute=-8.387562066e-01 lute=-2.359457121e-7 ua1=1.731809447e-09 lua1=-4.504218931e-16 ub1=-7.088737332e-19 lub1=3.852747156e-26 uc1=7.631824104e-11 luc1=-3.531650240e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.114 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.303289752e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.152585767e-8 k1=4.221882219e-02 lk1=2.165518251e-7 k2=1.272986658e-01 lk2=-6.830565219e-08 wk2=-2.220446049e-22 pk2=-8.326672685e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383648e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267778e-8 nfactor=4.152229107e+00 lnfactor=-5.540174069e-7 eta0=9.800711344e-01 leta0=-2.452271850e-7 etab=4.281583539e-02 letab=-2.173740306e-08 wetab=8.326672685e-23 petab=1.734723476e-30 u0=1.871952528e-02 lu0=3.764314976e-10 ua=-1.777587834e-09 lua=1.668975788e-16 ub=1.993952344e-18 lub=-2.057068089e-25 uc=1.245140400e-11 luc=2.005847147e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.384900615e+05 lvsat=-2.629607820e-02 wvsat=1.862645149e-15 a0=1.269019515e+00 la0=5.783543445e-8 ags=-9.392106230e-01 lags=5.481586371e-07 wags=1.776356839e-21 a1=0.0 a2=0.42385546 b0=-4.603925132e-17 lb0=1.152781418e-23 b1=1.027396975e-17 lb1=-2.572509561e-24 keta=6.904029211e-02 lketa=-3.810657865e-08 wketa=-1.110223025e-22 pketa=-8.326672685e-29 dwg=0.0 dwb=0.0 pclm=6.653835068e-01 lpclm=-1.068702608e-7 pdiblc1=-2.914152067e-01 lpdiblc1=1.623503586e-07 wpdiblc1=2.220446049e-22 ppdiblc1=2.220446049e-28 pdiblc2=-8.326311299e-03 lpdiblc2=4.189648227e-09 wpdiblc2=5.204170428e-24 ppdiblc2=-8.673617380e-31 pdiblcb=-8.590105794e-02 lpdiblcb=-4.355479349e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974521e+07 lpscbe1=1.776524482e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465818e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-06 wbeta0=-1.136868377e-19 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-08 wkt1=1.776356839e-21 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438220939e+03 lat=9.053815040e-3 ute=-1.301500893e+00 lute=-4.392435834e-9 ua1=1.688524505e-09 lua1=-4.287624978e-16 ub1=-1.973606354e-18 lub1=6.713882924e-25 wub1=6.162975822e-39 pub1=-1.540743956e-45 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=1.033975766e-31 puc1=1.809457590e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.115 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.724754252e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322497667e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232475895e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767208767e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665316856e-16 ags=1.250000000e+00 lags=5.707079254e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.562927813e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223410262e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387237549e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448285936e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435023e-25 ub1=7.077531678e-19 lub1=3.881565432e-34 uc1=1.471862500e-10 luc1=-5.619865082e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.116 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.993815894e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.882962214e-09 wvth0=9.255575520e-08 pvth0=-1.669622524e-14 k1=0.90707349 k2=-1.114045584e-01 lk2=-5.540854324e-09 wk2=-3.054881216e-09 pk2=5.510730774e-16 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585025681e-01 ldsub=2.298756365e-11 wdsub=7.026958387e-11 pdsub=-1.267600050e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.839084440e-19 cit=0.0 voff='-5.767390087e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.660198229e-08 wvoff=2.035235549e-07 pvoff=-3.671381760e-14 nfactor=-1.428319319e+01 lnfactor=2.980600330e-06 wnfactor=9.108104482e-06 pnfactor=-1.643020076e-12 eta0=1.783336336e-02 leta0=-3.216978204e-09 weta0=-9.830499004e-09 peta0=1.773333546e-15 etab=-0.043998 u0=-7.642541265e-02 lu0=1.844721445e-08 wu0=6.153667580e-08 pu0=-1.110066248e-14 ua=-6.409625481e-10 lua=-7.676553370e-17 wua=-2.595732714e-16 pua=4.682468201e-23 ub=2.506649802e-17 lub=-4.230263817e-24 wub=-1.282427509e-23 pub=2.313383808e-30 uc=3.478607631e-10 luc=-4.886012235e-17 wuc=-1.493584271e-16 puc=2.694291603e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.486150032e+06 lvsat=-5.846705881e-01 wvsat=-1.839120929e+00 pvsat=3.317608634e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000008e-02 lketa=1.268496419e-17 dwg=0.0 dwb=0.0 pclm=-3.426699911e-01 lpclm=9.415803752e-08 wpclm=2.775781595e-07 ppclm=-5.007260176e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.786314880e-24 alpha1=0.85 beta0=1.392897432e+01 lbeta0=-1.187702761e-8 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.918229421e-01 lkt1=4.693873204e-08 wkt1=1.416215050e-07 pkt1=-2.554724491e-14 kt2=-0.028878939 at=5.372048691e+04 lat=1.396238804e-11 ute=3.516368414e-01 lute=-3.007833360e-07 wute=-9.103751749e-07 pute=1.642234882e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.117 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.118 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-6 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 wub=-3.081487911e-39 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-7 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 wb0=1.499264860e-30 pb0=2.192028623e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-7 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+03 ppscbe1=7.629394531e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-8 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344737e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.119 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008797e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 wb0=-1.323488980e-29 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539119e-02 lketa=8.113189461e-08 wketa=2.775557562e-23 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=-8.881784197e-22 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 uc1=-7.151779256e-11 luc1=4.155336487e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.120 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155422e-01 leta0=-3.180932596e-7 etab=-1.395135872e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 b1=-5.828486835e-09 lb1=5.498972206e-14 pb1=5.293955920e-35 keta=4.904572511e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-6 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-8 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-01 wat=-4.656612873e-16 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 pua1=6.617444900e-36 ub1=-1.496090981e-18 lub1=3.294685946e-24 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.121 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-09 peta0=1.734723476e-30 etab=8.340779512e-02 letab=-1.678483982e-07 wetab=-1.040834086e-22 petab=-1.474514955e-28 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 ub=-4.679975144e-19 lub=1.932152691e-24 pub=-1.540743956e-45 uc=6.203139367e-11 luc=-2.248718272e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024581e-01 lags=1.548007492e-6 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 pb0=1.058791184e-34 b1=3.210308126e-08 lb1=-2.088824537e-14 keta=7.274507804e-02 lketa=-1.354760365e-07 wketa=5.551115123e-23 pketa=-2.775557562e-29 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-9 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=-2.117582368e-28 palpha0=7.411538288e-34 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-8 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-6 ua1=-1.595365930e-09 lua1=2.878054409e-15 wua1=8.271806126e-31 pua1=3.308722450e-36 ub1=9.725424449e-19 lub1=-1.643546140e-24 wub1=7.703719778e-40 pub1=7.703719778e-46 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.122 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.027376911e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.355915084e-08 wvth0=2.171702671e-08 pvth0=-2.172551806e-14 k1=6.334555289e-01 lk1=-7.929770217e-08 wk1=-3.737543608e-16 pk1=3.739017984e-22 k2=-7.088141908e-02 lk2=2.888185447e-08 wk2=-2.024543070e-09 pk2=2.025334666e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535300e-01 ldsub=5.036615542e-08 wdsub=-1.102380409e-16 pdsub=1.102806735e-22 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891544e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980655631e-09 wvoff=-4.547744403e-16 pvoff=4.549520760e-22 nfactor=2.048395165e+00 lnfactor=4.987221588e-07 wnfactor=-4.418680533e-15 pnfactor=4.420414257e-21 eta0=-4.853187011e-01 leta0=4.880407004e-07 weta0=2.522196618e-16 peta0=-2.523184786e-22 etab=-1.681904926e-01 letab=8.384826446e-08 wetab=5.067635200e-17 petab=-5.069611397e-23 u0=-8.682674873e-03 lu0=3.023079049e-08 wu0=1.650549363e-08 pu0=-1.651194728e-14 ua=-7.984359590e-10 lua=-3.230612086e-16 wua=-1.588468018e-24 pua=1.589090057e-30 ub=1.343841469e-18 lub=1.196052787e-25 wub=2.512008077e-30 pub=-2.512990274e-36 uc=2.655884663e-11 luc=1.299923409e-17 wuc=-5.681035088e-26 puc=5.683258136e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.653606010e+06 lvsat=1.737701185e+00 wvsat=7.844193757e-01 pvsat=-7.847260837e-7 a0=1.015255637e+00 la0=1.848165978e-07 wa0=2.747647443e-15 pa0=-2.748720362e-21 ags=2.344605288e+00 lags=-1.095033278e-06 wags=1.214111478e-14 pags=-1.214586121e-20 a1=0.0 a2=0.42385546 b0=1.610149328e-07 lb0=-8.057042354e-14 wb0=-2.890614282e-22 pb0=2.891745071e-28 b1=2.245477625e-08 lb1=-1.123616788e-14 wb1=6.450600586e-23 pb1=-6.453125803e-29 keta=-1.182861553e-01 lketa=5.562989013e-08 wketa=4.189208980e-16 pketa=-4.190846559e-22 dwg=0.0 dwb=0.0 pclm=1.289197297e+00 lpclm=-4.190210702e-07 wpclm=-3.209471799e-15 ppclm=3.210727684e-21 pdiblc1=6.759562110e-01 lpdiblc1=-3.217135918e-07 wpdiblc1=6.015863363e-16 ppdiblc1=-6.018225918e-22 pdiblc2=9.346473056e-03 lpdiblc2=-4.653654024e-09 wpdiblc2=-1.449775022e-17 ppdiblc2=1.450341930e-23 pdiblcb=9.429603766e-02 lpdiblcb=-9.452448410e-08 wpdiblcb=1.164782819e-16 ppdiblcb=-1.165240560e-22 drout=8.393443491e-01 ldrout=8.039059138e-08 wdrout=-4.043059221e-16 pdrout=4.044640178e-22 pscbe1=1.031079496e+09 lpscbe1=-2.972985438e+02 wpscbe1=4.655429840e-06 ppscbe1=-4.657251358e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266829e-06 lalpha0=-1.621900744e-12 walpha0=5.464514475e-21 palpha0=-5.466642221e-27 alpha1=0.85 beta0=1.690956682e+01 lbeta0=5.546499618e-07 wbeta0=-2.433097279e-14 pbeta0=2.434049406e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611033e-01 lkt1=-4.297596406e-09 wkt1=3.904521151e-17 pkt1=-3.906031054e-23 kt2=-1.752560649e-02 lkt2=-9.604001211e-09 wkt2=6.363909399e-18 pkt2=-6.366407401e-24 at=1.147614886e+05 lat=-5.209381936e-02 wat=4.835315049e-10 pat=-4.837205634e-16 ute=-8.387562047e-01 lute=-2.359457141e-07 wute=-9.994529648e-16 pute=9.998437633e-22 ua1=1.731809443e-09 lua1=-4.504218890e-16 wua1=2.070538952e-24 pua1=-2.071349589e-30 ub1=-7.088737341e-19 lub1=3.852747245e-26 wub1=4.542729478e-34 pub1=-4.544501334e-40 uc1=7.631824114e-11 luc1=-3.531650250e-17 wuc1=-5.031305396e-26 puc1=5.033259611e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.123 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='7.152868883e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.279855449e-08 wvth0=-4.343405341e-08 pvth0=1.087549607e-14 k1=4.221882073e-02 lk1=2.165518255e-07 wk1=7.475104979e-16 pk1=-1.871698352e-22 k2=1.193785690e-01 lk2=-6.632253122e-08 wk2=4.049086140e-09 pk2=-1.013854728e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522826e-01 ldsub=7.433550855e-08 wdsub=2.204743055e-16 pdsub=-5.520495172e-23 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383665e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267733e-08 wvoff=9.095488807e-16 pvoff=-2.277428246e-22 nfactor=4.152229090e+00 lnfactor=-5.540174026e-07 wnfactor=8.837375276e-15 pnfactor=-2.212797057e-21 eta0=9.800711353e-01 leta0=-2.452271852e-07 weta0=-5.044391571e-16 peta0=1.263069649e-22 etab=4.281583558e-02 letab=-2.173740311e-08 wetab=-1.013524195e-16 petab=2.537771729e-23 u0=8.328970391e-02 lu0=-1.579136010e-08 wu0=-3.301098726e-08 pu0=8.265654112e-15 ua=-1.777587840e-09 lua=1.668975804e-16 wua=3.176936035e-24 pua=-7.954764340e-31 ub=1.993962171e-18 lub=-2.057092695e-25 wub=-5.024016154e-30 pub=1.257968429e-36 uc=1.245140378e-11 luc=2.005847152e-17 wuc=1.136207018e-25 puc=-2.844958470e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.407171335e+06 lvsat=-7.946662508e-01 wvsat=-1.568838751e+00 pvsat=3.928231038e-7 a0=1.269019526e+00 la0=5.783543176e-08 wa0=-5.495294886e-15 pa0=1.375971337e-21 ags=-9.392105755e-01 lags=5.481586252e-07 wags=-2.428222823e-14 pags=6.080051018e-21 a1=0.0 a2=0.42385546 b0=-1.176859946e-15 lb0=2.946751388e-22 wb0=5.781230337e-22 pb0=-1.447568045e-28 b1=2.626242423e-16 lb1=-6.575874664e-23 wb1=-1.290120580e-22 pb1=3.230345822e-29 keta=6.904029375e-02 lketa=-3.810657906e-08 wketa=-8.378416849e-16 pketa=2.097880411e-22 dwg=0.0 dwb=0.0 pclm=6.653834942e-01 lpclm=-1.068702576e-07 wpclm=6.418945375e-15 ppclm=-1.607245892e-21 pdiblc1=-2.914152043e-01 lpdiblc1=1.623503581e-07 wpdiblc1=-1.203174227e-15 ppdiblc1=3.012642080e-22 pdiblc2=-8.326311356e-03 lpdiblc2=4.189648241e-09 wpdiblc2=2.899549437e-17 ppdiblc2=-7.260206433e-24 pdiblcb=-8.590105748e-02 lpdiblcb=-4.355479463e-09 wpdiblcb=-2.329567650e-16 ppdiblcb=5.833034056e-23 drout=1.497449936e+00 ldrout=-2.489195212e-07 wdrout=8.086118441e-16 pdrout=-2.024691526e-22 pscbe1=8.191976342e+07 lpscbe1=1.776524437e+02 wpscbe1=-9.310861588e-06 ppscbe1=2.331356525e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465840e-06 lalpha0=-1.943751740e-12 walpha0=-1.092902895e-20 palpha0=2.736529671e-27 alpha1=0.85 beta0=2.172178357e+01 lbeta0=-1.853339991e-06 wbeta0=4.866194558e-14 pbeta0=-1.218451473e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978344e-01 lkt1=1.903900409e-08 wkt1=-7.809042302e-17 pkt1=1.955302587e-23 kt2=-4.457052220e-02 lkt2=3.929031209e-09 wkt2=-1.272770778e-17 pkt2=3.186950703e-24 at=-7.438219047e+03 lat=9.053814566e-03 wat=-9.670630679e-10 pat=2.421438985e-16 ute=-1.301500897e+00 lute=-4.392434855e-09 wute=1.998913035e-15 pute=-5.005098558e-22 ua1=1.688524513e-09 lua1=-4.287624998e-16 wua1=-4.141077905e-24 pua1=1.036888269e-30 ub1=-1.973606352e-18 lub1=6.713882920e-25 wub1=-9.085458957e-34 pub1=2.274923858e-40 uc1=-1.359266153e-10 luc1=7.088891345e-17 wuc1=1.006258753e-25 puc1=-2.519584391e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.124 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.724931888e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322408849e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232475895e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767319789e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665281329e-16 ags=1.250000000e+00 lags=5.706368711e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.563016631e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223410262e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387428284e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448174913e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435540e-25 ub1=7.077531678e-19 lub1=3.881565432e-34 uc1=1.471862500e-10 luc1=-5.620278672e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.125 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.069683588e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.524722703e-09 wvth0=3.755288005e-08 pvth0=-6.774201585e-15 k1=0.90707349 k2=-4.183667196e-01 lk2=4.983235690e-08 wk2=1.538770680e-07 pk2=-2.775803817e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585032325e-01 ldsub=2.286771234e-11 wdsub=6.992991602e-11 pdsub=-1.261472748e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.839223218e-19 cit=0.0 voff='-5.767412486e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.660238635e-08 wvoff=2.035247001e-07 pvoff=-3.671402417e-14 nfactor=-1.428319340e+01 lnfactor=2.980600368e-06 wnfactor=9.108104589e-06 pnfactor=-1.643020095e-12 eta0=1.783336150e-02 leta0=-3.216977870e-09 weta0=-9.830498056e-09 peta0=1.773333375e-15 etab=-0.043998 u0=4.339052496e-01 lu0=-7.361184404e-08 wu0=-1.993657926e-07 pu0=3.596379470e-14 ua=-6.409392434e-10 lua=-7.676973766e-17 wua=-2.595851858e-16 pua=4.682683125e-23 ub=2.506644320e-17 lub=-4.230253928e-24 wub=-1.282424706e-23 pub=2.313378752e-30 uc=3.464485825e-10 luc=-4.860537769e-17 wuc=-1.486364611e-16 puc=2.681267986e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.723447900e+06 lvsat=3.550939925e-01 wvsat=8.242443374e-01 pvsat=-1.486862603e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000008e-02 lketa=1.268474215e-17 dwg=0.0 dwb=0.0 pclm=-3.426700025e-01 lpclm=9.415803956e-08 wpclm=2.775781653e-07 ppclm=-5.007260281e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.786209001e-24 alpha1=0.85 beta0=1.392897432e+01 lbeta0=-1.187702761e-8 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.918229625e-01 lkt1=4.693873572e-08 wkt1=1.416215154e-07 pkt1=-2.554724679e-14 kt2=-0.028878939 at=5.372048691e+04 lat=1.396285370e-11 ute=3.430292648e-01 lute=-2.992306067e-07 wute=-9.059746203e-07 pute=1.634296677e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.126 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.127 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-07 pk2=4.440892099e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-06 wnfactor=7.105427358e-21 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-7 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 wb0=7.496324301e-31 pb0=1.571643164e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-07 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+03 ppscbe1=3.814697266e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-08 wkt1=-4.440892099e-22 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344738e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 puc1=4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.128 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-07 pk2=1.110223025e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008798e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 pb0=-5.293955920e-35 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539119e-02 lketa=8.113189461e-08 wketa=-1.387778781e-23 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=-2.220446049e-22 ppclm=1.332267630e-27 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-08 ppdiblc2=-1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 wub1=1.540743956e-39 uc1=-7.151779256e-11 luc1=4.155336487e-16 wuc1=5.169878828e-32 puc1=-2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.129 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155422e-01 leta0=-3.180932596e-7 etab=-1.395135872e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 wb0=-1.323488980e-29 pb0=-2.646977960e-35 b1=-5.828486835e-09 lb1=5.498972206e-14 keta=4.904572512e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-6 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-8 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-1 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 ub1=-1.496090981e-18 lub1=3.294685946e-24 pub1=-3.081487911e-45 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.130 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-9 etab=8.340779513e-02 letab=-1.678483982e-07 wetab=-2.428612866e-23 petab=-4.163336342e-29 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 ub=-4.679975144e-19 lub=1.932152691e-24 pub=-1.540743956e-45 uc=6.203139367e-11 luc=-2.248718272e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024580e-01 lags=1.548007492e-06 pags=-8.881784197e-28 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 b1=3.210308126e-08 lb1=-2.088824537e-14 keta=7.274507804e-02 lketa=-1.354760365e-07 pketa=-5.551115123e-29 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-9 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=1.270549421e-27 palpha0=1.747005454e-33 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-8 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-6 ua1=-1.595365930e-09 lua1=2.878054409e-15 wua1=8.271806126e-31 ub1=9.725424449e-19 lub1=-1.643546140e-24 pub1=3.851859889e-46 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.131 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.469460990e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.933345747e-8 k1=6.334555281e-01 lk1=-7.929770141e-8 k2=-7.500269346e-02 lk2=3.300474027e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615565e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891554e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980654705e-9 nfactor=2.048395156e+00 lnfactor=4.987221678e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=9.020562075e-23 peta0=1.457167720e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.491684152e-02 lu0=-3.381863310e-9 ua=-7.984359622e-10 lua=-3.230612054e-16 ub=1.343846582e-18 lub=1.196001631e-25 uc=2.655884651e-11 luc=1.299923420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.679756133e+04 lvsat=1.402683848e-01 pvsat=-1.164153218e-22 a0=1.015255643e+00 la0=1.848165922e-7 ags=2.344605312e+00 lags=-1.095033303e-6 a1=0.0 a2=0.42385546 b0=1.610149322e-07 lb0=-8.057042295e-14 b1=2.245477639e-08 lb1=-1.123616801e-14 keta=-1.182861545e-01 lketa=5.562988928e-8 dwg=0.0 dwb=0.0 pclm=1.289197290e+00 lpclm=-4.190210637e-7 pdiblc1=6.759562122e-01 lpdiblc1=-3.217135930e-7 pdiblc2=9.346473027e-03 lpdiblc2=-4.653653994e-9 pdiblcb=9.429603790e-02 lpdiblcb=-9.452448434e-08 wpdiblcb=3.165870344e-23 ppdiblcb=-4.423544864e-29 drout=8.393443482e-01 ldrout=8.039059221e-8 pscbe1=1.031079505e+09 lpscbe1=-2.972985533e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266840e-06 lalpha0=-1.621900755e-12 alpha1=0.85 beta0=1.690956677e+01 lbeta0=5.546500114e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611032e-01 lkt1=-4.297596485e-9 kt2=-1.752560647e-02 lkt2=-9.604001224e-9 at=1.147614896e+05 lat=-5.209382035e-2 ute=-8.387562067e-01 lute=-2.359457120e-7 ua1=1.731809447e-09 lua1=-4.504218933e-16 ub1=-7.088737332e-19 lub1=3.852747153e-26 uc1=7.631824104e-11 luc1=-3.531650239e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.132 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.268700725e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.065977958e-8 k1=4.221882225e-02 lk1=2.165518251e-7 k2=1.276211178e-01 lk2=-6.838639125e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383647e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267780e-8 nfactor=4.152229108e+00 lnfactor=-5.540174071e-7 eta0=9.800711343e-01 leta0=-2.452271850e-7 etab=4.281583538e-02 letab=-2.173740306e-08 wetab=1.214306433e-23 petab=-8.673617380e-30 u0=1.609067113e-02 lu0=1.034672918e-9 ua=-1.777587834e-09 lua=1.668975787e-16 ub=1.993951944e-18 lub=-2.057067087e-25 uc=1.245140401e-11 luc=2.005847146e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.135544382e+05 lvsat=4.986677451e-3 a0=1.269019515e+00 la0=5.783543456e-8 ags=-9.392106249e-01 lags=5.481586376e-07 wags=-4.440892099e-22 pags=-3.330669074e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.904029204e-02 lketa=-3.810657863e-08 wketa=-1.387778781e-23 pketa=-1.040834086e-29 dwg=0.0 dwb=0.0 pclm=6.653835073e-01 lpclm=-1.068702609e-7 pdiblc1=-2.914152068e-01 lpdiblc1=1.623503587e-07 wpdiblc1=-1.665334537e-22 ppdiblc1=1.110223025e-28 pdiblc2=-8.326311297e-03 lpdiblc2=4.189648226e-09 ppdiblc2=3.523657061e-31 pdiblcb=-8.590105796e-02 lpdiblcb=-4.355479344e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974447e+07 lpscbe1=1.776524484e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465817e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-8 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438221016e+03 lat=9.053815059e-3 ute=-1.301500893e+00 lute=-4.392435874e-9 ua1=1.688524505e-09 lua1=-4.287624977e-16 ub1=-1.973606354e-18 lub1=6.713882925e-25 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=9.047287950e-32 puc1=2.261821987e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.133 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.724931888e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322408849e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232510589e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767264278e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665316856e-16 ags=1.250000000e+00 lags=5.706723982e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.562972222e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223438018e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416742362e-16 pscbe1=7.914198799e+08 lpscbe1=2.387523651e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448063891e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435023e-25 ub1=7.077531678e-19 lub1=3.881565432e-34 uc1=1.471862500e-10 luc1=-5.620278672e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.134 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.659102366e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.015730699e-08 wvth0=8.598154093e-09 pvth0=-1.551029615e-15 k1=0.90707349 k2=-2.070157960e-01 lk2=1.170655243e-08 wk2=5.005261758e-08 pk2=-9.029041738e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585044677e-01 ldsub=2.264489295e-11 wdsub=6.932313273e-11 pdsub=-1.250526924e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.839188524e-19 cit=0.0 voff='-5.767402513e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.660220644e-08 wvoff=2.035242101e-07 pvoff=-3.671393579e-14 nfactor=-1.428319270e+01 lnfactor=2.980600242e-06 wnfactor=9.108104246e-06 pnfactor=-1.643020033e-12 eta0=1.783333504e-02 leta0=-3.216973097e-09 weta0=-9.830485059e-09 peta0=1.773331030e-15 etab=-0.043998 u0=1.846997955e-01 lu0=-2.865742297e-08 wu0=-7.694560694e-08 pu0=1.388029498e-14 ua=-6.409159161e-10 lua=-7.677394570e-17 wua=-2.595966452e-16 pua=4.682889842e-23 ub=2.506645159e-17 lub=-4.230255441e-24 wub=-1.282425118e-23 pub=2.313379495e-30 uc=3.438160171e-10 luc=-4.813048659e-17 wuc=-1.473432344e-16 puc=2.657939340e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.377984282e+06 lvsat=2.927754650e-01 wvsat=6.545380988e-01 pvsat=-1.180727822e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000008e-02 lketa=1.268479766e-17 dwg=0.0 dwb=0.0 pclm=-3.426700067e-01 lpclm=9.415804032e-08 wpclm=2.775781673e-07 ppclm=-5.007260318e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.786261940e-24 alpha1=0.85 beta0=1.392897432e+01 lbeta0=-1.187702761e-8 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-4.918229539e-01 lkt1=4.693873418e-08 wkt1=1.416215112e-07 pkt1=-2.554724603e-14 kt2=-0.028878939 at=5.372048691e+04 lat=1.396285370e-11 ute=3.269831878e-01 lute=-2.963360388e-07 wute=-8.980921133e-07 pute=1.620077344e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.135 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.136 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-6 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-7 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 wb0=2.688336991e-30 pb0=-1.075334796e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-07 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+03 ppscbe1=-7.629394531e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-8 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344737e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.137 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008797e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 wb0=2.646977960e-29 pb0=-5.293955920e-35 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539119e-02 lketa=8.113189461e-8 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=-4.440892099e-22 ppclm=7.105427358e-27 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 uc1=-7.151779256e-11 luc1=4.155336487e-16 puc1=4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.138 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-06 wdsub=3.552713679e-21 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155422e-01 leta0=-3.180932596e-7 etab=-1.395135872e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 pb0=-1.058791184e-34 b1=-5.828486835e-09 lb1=5.498972206e-14 keta=4.904572512e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-6 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-8 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-1 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 ub1=-1.496090981e-18 lub1=3.294685946e-24 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.139 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-9 etab=8.340779512e-02 letab=-1.678483982e-07 wetab=-6.938893904e-24 petab=1.804112415e-28 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 ub=-4.679975144e-19 lub=1.932152691e-24 uc=6.203139367e-11 luc=-2.248718272e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024581e-01 lags=1.548007492e-06 pags=3.552713679e-27 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 b1=3.210308126e-08 lb1=-2.088824537e-14 keta=7.274507804e-02 lketa=-1.354760365e-07 wketa=8.326672685e-23 pketa=-1.110223025e-28 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-9 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=-3.176373552e-27 palpha0=-1.058791184e-33 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-8 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-6 ua1=-1.595365930e-09 lua1=2.878054409e-15 wua1=-1.654361225e-30 pua1=8.271806126e-37 ub1=9.725424449e-19 lub1=-1.643546140e-24 wub1=7.703719778e-40 pub1=7.703719778e-46 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.140 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.469460990e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.933345747e-8 k1=6.334555281e-01 lk1=-7.929770141e-8 k2=-7.500269346e-02 lk2=3.300474027e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615565e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891554e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980654705e-9 nfactor=2.048395156e+00 lnfactor=4.987221678e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=3.608224830e-22 peta0=-5.065392550e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.491684152e-02 lu0=-3.381863310e-09 wu0=1.110223025e-22 ua=-7.984359622e-10 lua=-3.230612054e-16 ub=1.343846582e-18 lub=1.196001631e-25 uc=2.655884651e-11 luc=1.299923420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.679756133e+04 lvsat=1.402683848e-01 pvsat=2.328306437e-22 a0=1.015255643e+00 la0=1.848165922e-7 ags=2.344605313e+00 lags=-1.095033303e-6 a1=0.0 a2=0.42385546 b0=1.610149322e-07 lb0=-8.057042295e-14 b1=2.245477639e-08 lb1=-1.123616801e-14 keta=-1.182861545e-01 lketa=5.562988928e-8 dwg=0.0 dwb=0.0 pclm=1.289197290e+00 lpclm=-4.190210637e-7 pdiblc1=6.759562122e-01 lpdiblc1=-3.217135930e-7 pdiblc2=9.346473027e-03 lpdiblc2=-4.653653994e-9 pdiblcb=9.429603790e-02 lpdiblcb=-9.452448434e-08 wpdiblcb=-4.857225733e-23 ppdiblcb=-7.459310947e-29 drout=8.393443482e-01 ldrout=8.039059221e-8 pscbe1=1.031079505e+09 lpscbe1=-2.972985533e+02 wpscbe1=3.814697266e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266840e-06 lalpha0=-1.621900755e-12 alpha1=0.85 beta0=1.690956677e+01 lbeta0=5.546500114e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611032e-01 lkt1=-4.297596485e-9 kt2=-1.752560647e-02 lkt2=-9.604001224e-9 at=1.147614896e+05 lat=-5.209382035e-2 ute=-8.387562067e-01 lute=-2.359457120e-7 ua1=1.731809447e-09 lua1=-4.504218933e-16 ub1=-7.088737332e-19 lub1=3.852747153e-26 uc1=7.631824104e-11 luc1=-3.531650239e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.141 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.268700725e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.065977958e-8 k1=4.221882225e-02 lk1=2.165518251e-7 k2=1.276211178e-01 lk2=-6.838639125e-08 wk2=-2.220446049e-22 pk2=-8.326672685e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-09 pcdscd=6.938893904e-30 cit=0.0 voff='-1.087383647e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267780e-8 nfactor=4.152229108e+00 lnfactor=-5.540174071e-07 wnfactor=1.421085472e-20 eta0=9.800711343e-01 leta0=-2.452271850e-7 etab=4.281583538e-02 letab=-2.173740306e-08 wetab=-3.816391647e-23 petab=-2.688821388e-29 u0=1.609067113e-02 lu0=1.034672918e-9 ua=-1.777587834e-09 lua=1.668975787e-16 ub=1.993951944e-18 lub=-2.057067087e-25 uc=1.245140401e-11 luc=2.005847146e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.135544382e+05 lvsat=4.986677451e-3 a0=1.269019515e+00 la0=5.783543456e-8 ags=-9.392106249e-01 lags=5.481586376e-07 wags=1.776356839e-21 pags=4.440892099e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.904029204e-02 lketa=-3.810657863e-08 wketa=-5.551115123e-23 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=6.653835073e-01 lpclm=-1.068702609e-7 pdiblc1=-2.914152068e-01 lpdiblc1=1.623503587e-07 ppdiblc1=1.110223025e-28 pdiblc2=-8.326311297e-03 lpdiblc2=4.189648226e-09 wpdiblc2=-1.105886216e-23 ppdiblc2=4.336808690e-30 pdiblcb=-8.590105796e-02 lpdiblcb=-4.355479344e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974447e+07 lpscbe1=1.776524484e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465817e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-8 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438221016e+03 lat=9.053815059e-3 ute=-1.301500893e+00 lute=-4.392435874e-9 ua1=1.688524505e-09 lua1=-4.287624977e-16 ub1=-1.973606354e-18 lub1=6.713882925e-25 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=-1.550963649e-31 puc1=2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.142 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.725109524e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322320031e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232545284e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767208767e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665316856e-16 ags=1.250000000e+00 lags=5.707079254e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.563105449e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223410262e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387237549e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448174913e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435023e-25 ub1=7.077531678e-19 lub1=3.881565432e-34 uc1=1.471862500e-10 luc1=-5.620692262e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.143 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='-5.669828605e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.022455117e-07 wvth0=5.772602320e-07 pvth0=-1.041325505e-13 k1=0.90707349 k2=2.666341992e-02 lk2=-3.044707500e-08 wk2=-5.773005131e-08 pk2=1.041398169e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.636924948e+00 ldsub=-3.929448039e-07 wdsub=-1.004709696e-06 pdsub=1.812405868e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.839084440e-19 cit=0.0 voff='4.807647755e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.610910810e-08 wvoff=-8.466750752e-08 pvoff=1.527325635e-14 nfactor=1.316115762e+01 lnfactor=-1.970113557e-06 wnfactor=-3.550382785e-06 pnfactor=6.404571009e-13 eta0=-1.234611579e-02 leta0=2.227128218e-09 weta0=4.089545203e-09 peta0=-7.377171488e-16 etab=-0.043998 u0=3.627160091e-01 lu0=-6.076994575e-08 wu0=-1.590541613e-07 pu0=2.869193922e-14 ua=-3.164017931e-09 lua=3.783709500e-16 wua=9.041639746e-16 pua=-1.631030435e-22 ub=-7.888276200e-18 lub=1.714480859e-24 wub=2.375853370e-24 pub=-4.285825653e-31 uc=-2.296160240e-10 luc=5.531149275e-17 wuc=1.171477071e-16 puc=-2.113239203e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.800393770e+06 lvsat=-6.413573303e-01 wvsat=-1.733947351e+00 pvsat=3.127884966e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.623720209e-01 lketa=1.506935942e-07 wketa=3.853086616e-07 pketa=-6.950621478e-14 dwg=0.0 dwb=0.0 pclm=8.779508459e-03 lpclm=3.075971083e-08 wpclm=1.154748901e-07 ppclm=-2.083063089e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.999997370e-08 lalpha0=4.745059301e-21 walpha0=1.213977276e-20 palpha0=-2.189905747e-27 alpha1=0.85 beta0=1.392897407e+01 lbeta0=-1.187698225e-08 wbeta0=1.159810381e-13 pbeta0=-2.092195928e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.847791130e-01 lkt1=-8.449211337e-09 wkt1=-4.051095459e-15 pkt1=7.307816574e-22 kt2=-0.028878939 at=5.372048974e+04 lat=-4.975781776e-10 wat=-1.307959668e-09 pat=2.359441714e-16 ute=-1.145176845e+00 lute=-3.077161832e-08 wute=-2.190700755e-07 pute=3.951826999e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.144 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.145 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.571856571e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.950165363e-7 k1=6.124668128e-01 lk1=-8.891992401e-7 k2=-4.676510727e-02 lk2=2.779806598e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016661769e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.322358477e-7 nfactor=4.254953535e+00 lnfactor=-8.267232321e-6 eta0=0.08 etab=-0.07 u0=1.873611106e-02 lu0=5.003675691e-8 ua=-1.234034189e-09 lua=3.757751243e-15 ub=1.359185733e-18 lub=-9.819338518e-25 uc=6.335039064e-11 luc=-2.962736048e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.391001388e+00 la0=-5.680388659e-7 ags=3.207921561e-01 lags=4.817662964e-7 a1=0.0 a2=0.42385546 b0=-1.749609710e-09 lb0=3.534820524e-14 wb0=8.271806126e-31 pb0=-2.316105715e-35 b1=1.181213187e-08 lb1=-2.668315903e-14 keta=-2.654640868e-03 lketa=-3.783992239e-8 dwg=0.0 dwb=0.0 pclm=-9.792970000e-03 lpclm=5.333698272e-07 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=5.504140665e-04 lpdiblc2=8.198428147e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.501413581e+07 lpscbe1=6.000400022e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832065116e-01 lkt1=-6.347100943e-8 kt2=-3.548263051e-02 lkt2=1.192963224e-7 at=1.983344738e+05 lat=-4.666985988e-1 ute=-1.015595122e+00 lute=-1.996136578e-6 ua1=1.029595533e-09 lua1=1.828125083e-15 ub1=-3.821008428e-19 lub1=-3.747456406e-24 uc1=6.941809319e-11 luc1=-7.120085432e-16 wuc1=-1.033975766e-31 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.146 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.046357902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.153969181e-7 k1=4.365554697e-01 lk1=5.181602866e-7 k2=1.942866573e-02 lk2=-2.515954060e-07 pk2=-1.110223025e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179970607e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.582391992e-9 nfactor=3.716618783e+00 lnfactor=-3.960343819e-6 eta0=0.08 etab=-0.07 u0=2.323312824e-02 lu0=1.405886115e-8 ua=-9.715491229e-10 lua=1.657768083e-15 ub=1.411757135e-18 lub=-1.402525622e-24 uc=9.497355943e-12 luc=1.345717293e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.410008797e+00 la0=-7.201055734e-7 ags=3.608480294e-01 lags=1.613036485e-7 a1=0.0 a2=0.42385546 b0=1.224923641e-08 lb0=-7.664803724e-14 wb0=6.617444900e-30 pb0=-5.293955920e-35 b1=9.036254672e-09 lb1=-4.475056080e-15 keta=-1.752539119e-02 lketa=8.113189461e-8 dwg=0.0 dwb=0.0 pclm=-6.991438936e-01 lpclm=6.048446752e-06 wpclm=2.220446049e-22 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.662990699e-03 lpdiblc2=2.590653171e-08 ppdiblc2=-1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.387919311e+08 lpscbe1=2.896723884e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862395210e-01 lkt1=-3.920574789e-8 kt2=-9.729417308e-03 lkt2=-8.673945272e-8 at=140000.0 ute=-1.230796647e+00 lute=-2.744402352e-7 ua1=1.517475351e-09 lua1=-2.075104227e-15 ub1=-1.028537400e-18 lub1=1.424288813e-24 uc1=-7.151779256e-11 luc1=4.155336487e-16 puc1=-2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.147 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.399336610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.580836658e-8 k1=5.590655484e-01 lk1=2.807207026e-8 k2=-4.343904111e-02 lk2=-9.999731753e-11 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.600586500e-01 ldsub=-1.200351923e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374705590e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.631921551e-8 nfactor=2.156847829e+00 lnfactor=2.279349867e-6 eta0=1.595155422e-01 leta0=-3.180932596e-7 etab=-1.395135872e-01 letab=2.780815288e-7 u0=2.768018230e-02 lu0=-3.731093894e-9 ua=-8.165774186e-10 lua=1.037820672e-15 wua=-1.654361225e-30 ub=1.624540119e-18 lub=-2.253740759e-24 uc=3.548250384e-11 luc=3.062097755e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.615275307e+00 la0=-1.541251869e-6 ags=3.258752828e-01 lags=3.012083092e-7 a1=0.0 a2=0.42385546 b0=-3.402409959e-08 lb0=1.084633996e-13 pb0=-5.293955920e-35 b1=-5.828486835e-09 lb1=5.498972206e-14 keta=4.904572511e-04 lketa=9.061456666e-9 dwg=0.0 dwb=0.0 pclm=1.120060054e+00 lpclm=-1.229080346e-6 pdiblc1=0.39 pdiblc2=2.445481039e-03 lpdiblc2=9.471038349e-9 pdiblcb=-3.750244375e-02 lpdiblcb=5.001466346e-8 drout=0.56 pscbe1=6.223885402e+08 lpscbe1=3.552923657e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.582526140e-01 lkt1=-1.511643188e-7 kt2=-1.455640634e-02 lkt2=-6.742960922e-8 at=1.706359882e+05 lat=-1.225559313e-1 ute=-8.683157395e-01 lute=-1.724505596e-6 ua1=2.154345875e-09 lua1=-4.622835337e-15 pua1=6.617444900e-36 ub1=-1.496090981e-18 lub1=3.294685946e-24 pub1=3.081487911e-45 uc1=8.123422561e-12 luc1=9.693764848e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.148 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.877766572e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.852603452e-8 k1=5.920162538e-01 lk1=-3.784222434e-8 k2=-4.496778497e-02 lk2=2.958088128e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.395669898e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.073724848e-8 nfactor=4.045970607e+00 lnfactor=-1.499634334e-6 eta0=-1.532044219e-03 leta0=4.064882967e-09 peta0=-1.734723476e-30 etab=8.340779513e-02 letab=-1.678483982e-07 wetab=-4.683753385e-23 petab=8.673617380e-30 u0=3.009537297e-02 lu0=-8.562419569e-9 ua=5.261559085e-10 lua=-1.648170992e-15 pua=8.271806126e-37 ub=-4.679975144e-19 lub=1.932152691e-24 uc=6.203139367e-11 luc=-2.248718272e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.658266434e+04 lvsat=6.836007490e-3 a0=4.894611168e-01 la0=7.108167039e-7 ags=-2.974024580e-01 lags=1.548007492e-6 a1=0.0 a2=0.42385546 b0=-4.010556909e-08 lb0=1.206287165e-13 pb0=5.293955920e-35 b1=3.210308126e-08 lb1=-2.088824537e-14 keta=7.274507804e-02 lketa=-1.354760365e-07 wketa=2.775557562e-23 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=1.407974023e-01 lpclm=7.298278489e-7 pdiblc1=4.256455720e-01 lpdiblc1=-7.130508136e-8 pdiblc2=9.666483106e-03 lpdiblc2=-4.973789197e-9 pdiblcb=-2.481331081e-02 lpdiblcb=2.463143613e-8 drout=2.001558359e-01 ldrout=7.198290272e-7 pscbe1=8.661286962e+08 lpscbe1=-1.322832487e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.462146590e-06 lalpha0=1.098644061e-11 walpha0=-1.588186776e-27 palpha0=6.352747104e-33 alpha1=0.85 beta0=1.025459084e+01 lbeta0=7.212228043e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.930061127e-01 lkt1=1.183953672e-7 kt2=-6.941165326e-02 lkt2=4.230233301e-08 wkt2=1.110223025e-22 at=1.560702227e+05 lat=-9.341870509e-2 ute=-2.386446714e+00 lute=1.312349942e-6 ua1=-1.595365930e-09 lua1=2.878054409e-15 wua1=4.135903063e-31 pua1=-4.135903063e-37 ub1=9.725424449e-19 lub1=-1.643546140e-24 pub1=-7.703719778e-46 uc1=7.215609079e-11 luc1=-3.115272474e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.149 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.469460990e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.933345747e-8 k1=6.334555281e-01 lk1=-7.929770141e-8 k2=-7.500269346e-02 lk2=3.300474027e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.096535298e-01 ldsub=5.036615565e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.256891554e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.980654705e-9 nfactor=2.048395156e+00 lnfactor=4.987221678e-7 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-2.706168623e-22 peta0=-3.469446952e-28 etab=-1.681904925e-01 letab=8.384826436e-8 u0=2.491684152e-02 lu0=-3.381863310e-9 ua=-7.984359622e-10 lua=-3.230612054e-16 ub=1.343846582e-18 lub=1.196001631e-25 uc=2.655884651e-11 luc=1.299923420e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.679756133e+04 lvsat=1.402683848e-01 pvsat=-1.164153218e-22 a0=1.015255643e+00 la0=1.848165922e-7 ags=2.344605313e+00 lags=-1.095033303e-6 a1=0.0 a2=0.42385546 b0=1.610149322e-07 lb0=-8.057042295e-14 b1=2.245477639e-08 lb1=-1.123616801e-14 keta=-1.182861545e-01 lketa=5.562988928e-8 dwg=0.0 dwb=0.0 pclm=1.289197290e+00 lpclm=-4.190210637e-7 pdiblc1=6.759562122e-01 lpdiblc1=-3.217135930e-7 pdiblc2=9.346473027e-03 lpdiblc2=-4.653653994e-9 pdiblcb=9.429603790e-02 lpdiblcb=-9.452448434e-08 wpdiblcb=4.466912951e-23 ppdiblcb=4.423544864e-29 drout=8.393443482e-01 ldrout=8.039059221e-8 pscbe1=1.031079505e+09 lpscbe1=-2.972985533e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.141266840e-06 lalpha0=-1.621900755e-12 alpha1=0.85 beta0=1.690956677e+01 lbeta0=5.546500114e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.703611032e-01 lkt1=-4.297596485e-9 kt2=-1.752560647e-02 lkt2=-9.604001224e-9 at=1.147614896e+05 lat=-5.209382035e-2 ute=-8.387562067e-01 lute=-2.359457120e-7 ua1=1.731809447e-09 lua1=-4.504218933e-16 ub1=-7.088737332e-19 lub1=3.852747153e-26 uc1=7.631824104e-11 luc1=-3.531650239e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.150 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.268700725e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.065977958e-8 k1=4.221882225e-02 lk1=2.165518251e-7 k2=1.276211178e-01 lk2=-6.838639125e-08 wk2=2.775557562e-23 pk2=6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.617522830e-01 ldsub=7.433550844e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-9 cit=0.0 voff='-1.087383647e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.746267780e-8 nfactor=4.152229108e+00 lnfactor=-5.540174071e-07 wnfactor=-7.105427358e-21 eta0=9.800711343e-01 leta0=-2.452271850e-7 etab=4.281583538e-02 letab=-2.173740306e-08 wetab=-1.908195824e-23 petab=9.974659987e-30 u0=1.609067113e-02 lu0=1.034672918e-9 ua=-1.777587834e-09 lua=1.668975787e-16 ub=1.993951944e-18 lub=-2.057067087e-25 uc=1.245140401e-11 luc=2.005847146e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.135544382e+05 lvsat=4.986677451e-3 a0=1.269019515e+00 la0=5.783543456e-8 ags=-9.392106249e-01 lags=5.481586376e-07 pags=-3.330669074e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.904029204e-02 lketa=-3.810657863e-08 wketa=-2.775557562e-23 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=6.653835073e-01 lpclm=-1.068702609e-7 pdiblc1=-2.914152068e-01 lpdiblc1=1.623503587e-07 wpdiblc1=-2.220446049e-22 ppdiblc1=2.775557562e-29 pdiblc2=-8.326311297e-03 lpdiblc2=4.189648226e-09 wpdiblc2=3.794707604e-24 ppdiblc2=-2.059984128e-30 pdiblcb=-8.590105796e-02 lpdiblcb=-4.355479344e-9 drout=1.497449937e+00 ldrout=-2.489195216e-7 pscbe1=8.191974447e+07 lpscbe1=1.776524484e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.784465817e-06 lalpha0=-1.943751735e-12 alpha1=0.85 beta0=2.172178367e+01 lbeta0=-1.853340015e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.169978345e-01 lkt1=1.903900413e-8 kt2=-4.457052223e-02 lkt2=3.929031215e-9 at=-7.438221016e+03 lat=9.053815059e-03 pat=7.275957614e-24 ute=-1.301500893e+00 lute=-4.392435874e-9 ua1=1.688524505e-09 lua1=-4.287624977e-16 ub1=-1.973606354e-18 lub1=6.713882925e-25 wub1=1.540743956e-39 pub1=-3.851859889e-46 uc1=-1.359266151e-10 luc1=7.088891340e-17 wuc1=1.292469707e-32 puc1=-4.523643975e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.151 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.190848321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.328674550e-9 k1=9.070734895e-01 lk1=8.724931888e-17 k2=-1.541996849e-01 lk2=2.179001335e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.322408849e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999995e-03 lcdscd=9.232545284e-19 cit=0.0 voff='-1.036177348e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483744e-8 nfactor=1.166036626e+00 lnfactor=1.936983146e-7 eta0=2.482948249e-03 leta0=-4.479014728e-10 etab=-4.399800002e-02 letab=3.767097745e-18 u0=5.755347348e-03 lu0=3.622544975e-9 ua=-1.225785826e-09 lua=2.873132216e-17 ub=2.934407110e-20 lub=2.862134211e-25 uc=1.326480344e-10 luc=-1.003768301e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.037040644e+05 lvsat=7.453122379e-3 a0=1.499999999e+00 la0=2.665352383e-16 ags=1.250000000e+00 lags=5.706368711e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.278421980e-01 lketa=3.623012494e-8 dwg=0.0 dwb=0.0 pclm=3.913189391e-01 lpclm=-3.824695960e-8 pdiblc1=3.569721503e-01 lpdiblc1=-4.562927813e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223451895e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622657729e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387619019e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.691922970e-11 lalpha0=5.420193807e-15 alpha1=0.85 beta0=1.549735057e+01 lbeta0=-2.947979878e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.650385764e-01 lkt1=6.028873541e-9 kt2=-2.887893901e-02 lkt2=1.448174913e-18 at=-3.570487010e+04 lat=1.613152959e-2 ute=-1.327504733e+00 lute=2.118691750e-9 ua1=-2.384733751e-11 lua1=2.732435540e-25 ub1=7.077531678e-19 lub1=3.881550025e-34 uc1=1.471862500e-10 luc1=-5.620278672e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.152 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.903107479e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.151926038e-08 wvth0=1.001649495e-07 pvth0=-1.806885541e-14 k1=0.90707349 k2=-7.388582768e-02 lk2=-1.230889567e-08 wk2=-1.235800773e-08 pk2=2.229273372e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.623230066e+00 ldsub=-3.904743706e-07 wdsub=-9.985299903e-07 pdsub=1.801258235e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.839223218e-19 cit=0.0 voff='4.807716289e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.610923172e-08 wvoff=-8.466781677e-08 pvoff=1.527331213e-14 nfactor=1.316115444e+01 lnfactor=-1.970112984e-06 wnfactor=-3.550381351e-06 pnfactor=6.404568422e-13 eta0=-1.234617400e-02 leta0=2.227138719e-09 weta0=4.089571470e-09 peta0=-7.377218871e-16 etab=-0.043998 u0=-1.727194897e-01 lu0=3.581779930e-08 wu0=8.255682400e-08 pu0=-1.489250804e-14 ua=-3.163917149e-09 lua=3.783527697e-16 wua=9.041184973e-16 pua=-1.630948399e-22 ub=-7.888225705e-18 lub=1.714471751e-24 wub=2.375830584e-24 pub=-4.285784549e-31 uc=-2.280192365e-10 luc=5.502344665e-17 wuc=1.164271695e-16 puc=-2.100241353e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.667891792e+06 lvsat=-2.566731660e-01 wvsat=-7.716728934e-01 pvsat=1.392028449e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.623738877e-01 lketa=1.506939310e-07 wketa=3.853095040e-07 pketa=-6.950636674e-14 dwg=0.0 dwb=0.0 pclm=8.779510267e-03 lpclm=3.075971051e-08 wpclm=1.154748892e-07 ppclm=-2.083063074e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000013e-08 lalpha0=-2.200041026e-23 walpha0=2.151338749e-22 palpha0=-3.880819091e-29 alpha1=0.85 beta0=1.392897433e+01 lbeta0=-1.187702860e-08 wbeta0=3.899458534e-17 pbeta0=-7.034373084e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.847791218e-01 lkt1=-8.449209750e-09 wkt1=-8.004086283e-17 pkt1=1.443867248e-23 kt2=-0.028878939 at=5.372048690e+04 lat=1.514214091e-11 wat=-2.540741116e-11 pat=4.583213013e-18 ute=-1.148162955e+00 lute=-3.023295087e-08 wute=-2.177226170e-07 pute=3.927520060e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.153 nmos lmin=2.0e-05 lmax=0.0001 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.154 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.320325602e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.980883080e-07 wvth0=1.084707179e-08 pvth0=-2.169456770e-13 k1=7.973854253e-01 lk1=-4.587643792e-06 wk1=-7.974467227e-08 pk1=1.594924625e-12 k2=-1.252532858e-01 lk2=1.847774918e-06 wk2=3.384739907e-08 pk2=-6.769612157e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.014176007e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.372074678e-07 wvoff=-1.071964741e-10 pvoff=2.143971395e-15 nfactor=4.761557726e+00 lnfactor=-1.839951422e-05 wnfactor=-2.184690046e-07 pnfactor=4.369465513e-12 eta0=0.08 etab=-0.07 u0=1.459715041e-02 lu0=1.328175884e-07 wu0=1.784893672e-09 pu0=-3.569857133e-14 ua=-1.564392659e-09 lua=1.036504982e-14 wua=1.424644474e-16 pua=-2.849344651e-21 ub=1.375770726e-18 lub=-1.313640204e-24 wub=-7.152145703e-27 pub=1.430457106e-31 uc=6.331284804e-11 luc=-2.955227382e-16 wuc=1.618994367e-20 puc=-3.238052036e-25 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.099494181e+00 la0=5.262219248e-06 wa0=1.257101508e-07 pa0=-2.514252169e-12 ags=3.188708586e-01 lags=5.201929976e-07 wags=8.285441760e-10 pags=-1.657120748e-14 a1=0.0 a2=0.42385546 b0=3.109640648e-08 lb0=-6.215849614e-13 wb0=-1.416458172e-14 pb0=2.832971727e-19 b1=1.155750474e-08 lb1=-2.159051690e-14 wb1=1.098059121e-16 pb1=-2.196161175e-21 keta=-4.953131026e-03 lketa=8.130779465e-09 wketa=9.912054924e-10 pketa=-1.982449741e-14 dwg=0.0 dwb=0.0 pclm=4.907381865e-02 lpclm=-6.439889628e-07 wpclm=-2.538583167e-08 ppclm=5.077265593e-13 pdiblc1=0.39 pdiblc2=2.897970408e-03 lpdiblc2=-3.875361657e-08 wpdiblc2=-1.012364892e-09 ppdiblc2=2.024769367e-14 pdiblcb=-0.025 drout=0.56 pscbe1=-1.015746162e+08 lpscbe1=6.531620015e+03 wpscbe1=1.145399468e+01 ppscbe1=-2.290843722e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.988418981e-01 lkt1=2.492428348e-07 wkt1=6.742635363e-09 pkt1=-1.348553436e-13 kt2=-5.872724513e-02 lkt2=5.841977034e-07 wkt2=1.002405410e-08 pkt2=-2.004850013e-13 at=2.314602927e+05 lat=-1.129227930e+00 wat=-1.428524441e-02 pat=2.857104738e-7 ute=-6.567320837e-01 lute=-9.173537665e-06 wute=-1.547568145e-07 pute=3.095196800e-12 ua1=1.538408112e-09 lua1=-8.348325443e-15 wua1=-2.194213542e-16 pua1=4.388512878e-21 ub1=-8.279522819e-19 lub1=5.169746705e-24 wub1=1.922698663e-25 pub1=-3.845472504e-30 uc1=1.563015821e-10 luc1=-2.449712292e-15 wuc1=-3.746780951e-17 puc1=7.493708401e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.155 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.240328550e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=2.620499773e-07 wvth0=-8.364829033e-09 pvth0=-6.324295855e-14 k1=-1.294343125e-01 lk1=2.827276497e-06 wk1=2.440785656e-07 pk1=-9.957878927e-13 k2=2.626508355e-01 lk2=-1.255609722e-06 wk2=-1.048876149e-07 pk2=4.329731418e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.134533789e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.177895088e-07 wvoff=-1.149334223e-08 pvoff=9.323758946e-14 nfactor=3.129908078e+00 lnfactor=-5.345679068e-06 wnfactor=2.530142979e-07 pnfactor=5.974147433e-13 eta0=0.08 etab=-0.07 u0=3.107511104e-02 lu0=9.874604179e-10 wu0=-3.381792347e-09 pu0=5.636936993e-15 ua=-1.281906144e-10 lua=-1.125128097e-15 wua=-3.636916099e-16 pua=1.200101714e-21 ub=1.044011878e-18 lub=1.340560297e-24 wub=1.585871998e-25 pub=-1.182933858e-30 uc=-6.703696932e-11 luc=7.473267675e-16 wuc=3.300481550e-17 puc=-2.642457082e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.085765790e+00 la0=-2.628339256e-06 wa0=-2.914147971e-07 pa0=8.229105099e-13 ags=2.088259352e-01 lags=1.400595412e-06 wags=6.555831194e-08 pags=-5.344346589e-13 a1=0.0 a2=0.42385546 b0=-1.724569221e-07 lb0=1.006921257e-12 wb0=7.965305323e-14 pb0=-4.672805896e-19 b1=1.583926798e-08 lb1=-5.584629702e-14 wb1=-2.933745067e-15 pb1=2.215343668e-20 keta=-1.162208748e-02 lketa=6.148503865e-08 wketa=-2.545752497e-09 pketa=8.472549458e-15 dwg=0.0 dwb=0.0 pclm=-1.862544379e+00 lpclm=1.464970406e-05 wpclm=5.017071523e-07 ppclm=-3.709223406e-12 pdiblc1=0.39 pdiblc2=-3.626762360e-03 lpdiblc2=1.344679674e-08 wpdiblc2=8.468608185e-10 ppdiblc2=5.373161029e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.012635248e+09 lpscbe1=-2.382494556e+03 wpscbe1=-1.612169397e+02 ppscbe1=1.152350617e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.981676911e-01 lkt1=2.438489151e-07 wkt1=5.143927916e-09 pkt1=-1.220650590e-13 kt2=1.930287702e-02 lkt2=-4.007378353e-08 wkt2=-1.251994467e-08 pkt2=-2.012419651e-14 at=4.062254316e+04 lat=3.975486839e-01 wat=4.285573324e-02 pat=-1.714396896e-7 ute=-2.641310337e+00 lute=6.703864330e-06 wute=6.082727446e-07 pute=-3.009338017e-12 ua1=-1.401076708e-09 lua1=1.516870245e-14 wua1=1.258602227e-15 pua1=-7.436253681e-21 ub1=1.170164665e-18 lub1=-1.081597013e-23 wub1=-9.481726761e-25 pub1=5.278513748e-30 uc1=-2.680313861e-10 luc1=9.451173677e-16 wuc1=8.474491512e-17 puc1=-2.283787421e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.156 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.445790611e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.201819806e-07 wvth0=-4.512749163e-08 pvth0=8.382206606e-14 k1=6.835303979e-01 lk1=-4.249002143e-07 wk1=-5.367447065e-08 pk1=1.953406739e-13 k2=-1.126863885e-01 lk2=2.458859307e-07 wk2=2.986236459e-08 pk2=-1.060794636e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.853978923e+00 ldsub=-5.176421639e-06 wdsub=-4.286201666e-07 pdsub=1.714648257e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.231492810e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.094777992e-07 wvoff=3.694826345e-08 pvoff=-1.005477739e-13 nfactor=-3.842277725e-01 lnfactor=8.712238363e-06 wnfactor=1.095818525e-06 pnfactor=-2.774131701e-12 eta0=4.229044147e-01 leta0=-1.371751734e-06 weta0=-1.135843441e-07 peta0=4.543817880e-13 etab=-3.697717839e-01 letab=1.199204346e-06 wetab=9.929700525e-08 petab=-3.972268461e-13 u0=3.007463586e-02 lu0=4.989752351e-09 wu0=-1.032588939e-09 pu0=-3.760795176e-15 ua=-1.828633708e-09 lua=5.677309151e-15 wua=4.364411784e-16 pua=-2.000742291e-21 ub=3.857916205e-18 lub=-9.916157245e-24 wub=-9.631255698e-25 pub=3.304355810e-30 uc=1.711011944e-10 luc=-2.053189994e-16 wuc=-5.848447536e-17 puc=1.017472276e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.052885953e+05 lvsat=-9.012424691e-01 wvsat=-9.715390442e-02 pvsat=3.886536049e-7 a0=4.183526438e+00 la0=-1.102020207e-05 wa0=-1.107537755e-06 pa0=4.087721444e-12 ags=-4.790271487e-02 lags=2.427610394e-06 wags=1.611887713e-07 pags=-9.169938877e-13 a1=0.0 a2=0.42385546 b0=-2.118161744e-07 lb0=1.164373655e-12 wb0=7.667140991e-14 pb0=-4.553528505e-19 b1=-1.609118966e-08 lb1=7.188801835e-14 wb1=4.425708490e-15 pb1=-7.287255091e-21 keta=4.522930502e-02 lketa=-1.659427602e-07 wketa=-1.929327019e-08 pketa=7.546916851e-14 dwg=0.0 dwb=0.0 pclm=7.373348468e+00 lpclm=-2.229747856e-05 wpclm=-2.696680602e-06 ppclm=9.085578183e-12 pdiblc1=0.39 pdiblc2=1.294534317e-02 lpdiblc2=-5.284810506e-08 wpdiblc2=-4.527981544e-09 ppdiblc2=2.687463204e-14 pdiblcb=-7.891578848e-02 lpdiblcb=2.156842350e-07 wpdiblcb=1.785917361e-08 ppdiblcb=-7.144367736e-14 drout=0.56 pscbe1=3.406478843e+07 lpscbe1=1.532169904e+03 wpscbe1=2.537099114e+02 ppscbe1=-5.075190233e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.014566265e-01 lkt1=-5.430722572e-07 wkt1=-6.761701523e-08 pkt1=1.690071632e-13 kt2=1.258951814e-01 lkt2=-4.664846787e-07 wkt2=-6.056862361e-08 pkt2=1.720893063e-13 at=2.721152481e+05 lat=-5.285126494e-01 wat=-4.376211901e-02 pat=1.750655870e-7 ute=1.607143079e+00 lute=-1.029161048e-05 wute=-1.067521812e-06 pute=3.694495444e-12 ua1=1.040453967e-08 lua1=-3.205837906e-14 wua1=-3.557830073e-15 pua1=1.183135875e-20 ub1=-6.673684046e-18 lub1=2.056249165e-23 wub1=2.232795589e-24 pub1=-7.446603069e-30 uc1=-1.577791545e-10 luc1=5.040653323e-16 wuc1=7.154415912e-17 puc1=-1.755705566e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.157 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.431429608e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.827689815e-07 wvth0=1.924792447e-08 pvth0=-4.495393693e-14 k1=4.921872138e-01 lk1=-4.213903081e-08 wk1=4.305047489e-08 pk1=1.852963413e-15 k2=1.757876805e-02 lk2=-1.469531614e-08 wk2=-2.697270062e-08 pk2=7.612889364e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.727840547e+00 ldsub=1.988617793e-06 wdsub=8.572403331e-07 pdsub=-8.575755141e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='4.784674676e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.326202159e-07 wvoff=-4.821434154e-08 pvoff=6.981073462e-14 nfactor=6.677944157e+00 lnfactor=-5.414866805e-06 wnfactor=-1.135017538e-06 pnfactor=1.688412681e-12 eta0=-5.283097891e-01 leta0=5.310485980e-07 weta0=2.271686883e-07 peta0=-2.272575112e-13 etab=8.224833688e-01 letab=-1.185772131e-06 wetab=-3.187204285e-07 petab=4.389714663e-13 u0=3.502585990e-02 lu0=-4.914631665e-09 wu0=-2.126233044e-09 pu0=-1.573079351e-15 ua=2.836438992e-09 lua=-3.654660293e-15 wua=-9.962910976e-16 pua=8.652824595e-22 ub=-3.858297774e-18 lub=5.519287752e-24 wub=1.462039865e-24 pub=-1.546923298e-30 uc=1.072832056e-10 luc=-7.765806901e-17 wuc=-1.951448189e-17 puc=2.379200335e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.719752226e+04 lvsat=-1.561245919e-01 wvsat=6.200405523e-02 pvsat=7.027545479e-8 a0=-2.857868091e+00 la0=3.065340170e-06 wa0=1.443508942e-06 pa0=-1.015369409e-12 ags=-2.390581297e+00 lags=7.113883545e-06 wags=9.026666287e-07 pags=-2.400239521e-12 a1=0.0 a2=0.42385546 b0=-6.644237705e-07 lb0=2.069765817e-12 wb0=2.692322298e-13 pb0=-8.405497815e-19 b1=4.611417868e-08 lb1=-5.254704063e-14 wb1=-6.042173676e-15 pb1=1.365260218e-20 keta=2.538969015e-01 lketa=-5.833595423e-07 wketa=-7.812027466e-08 pketa=1.931461788e-13 dwg=0.0 dwb=0.0 pclm=-7.871617123e+00 lpclm=8.198413405e-06 wpclm=3.455289665e-06 ppclm=-3.220767772e-12 pdiblc1=1.204491738e+00 lpdiblc1=-1.629301943e-06 wpdiblc1=-3.358711784e-07 ppdiblc1=6.718736825e-13 pdiblc2=-2.785900151e-02 lpdiblc2=2.877653880e-08 wpdiblc2=1.618256504e-08 ppdiblc2=-1.455455895e-14 pdiblcb=-2.419491782e-02 lpdiblcb=1.062210978e-07 wpdiblcb=-2.666770330e-10 ppdiblcb=-3.518488888e-14 drout=-6.795686010e-01 ldrout=2.479621873e-06 wdrout=3.793741256e-07 pdrout=-7.588965865e-13 pscbe1=1.085174712e+09 lpscbe1=-5.704609276e+02 wpscbe1=-9.446184199e+01 ppscbe1=1.889606186e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.365444280e-05 lalpha0=4.737814621e-11 walpha0=7.845282201e-12 palpha0=-1.569363191e-17 alpha1=0.85 beta0=-1.688038587e+00 lbeta0=3.110215646e-05 wbeta0=5.150163398e-06 pbeta0=-1.030234051e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-5.419069890e-01 lkt1=3.380006838e-07 wkt1=6.421231169e-08 pkt1=-9.470303594e-14 kt2=-1.852981043e-01 lkt2=1.560235693e-07 wkt2=4.997510492e-08 pkt2=-4.904137338e-14 at=1.761643980e+05 lat=-3.365734324e-01 wat=-8.665452366e-03 pat=1.048585309e-7 ute=-4.823701124e+00 lute=2.572592387e-06 wute=1.051046466e-06 pute=-5.434694725e-13 ua1=-9.502575809e-09 lua1=7.763635583e-15 wua1=3.409921003e-15 pua1=-2.106867797e-21 ub1=5.588457835e-18 lub1=-3.966586605e-24 wub1=-1.990576585e-24 pub1=1.001792616e-30 uc1=1.691066311e-10 luc1=-1.498340511e-16 wuc1=-4.180914489e-17 puc1=5.118037253e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.158 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.225180840e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.323722629e-09 wvth0=-3.258981398e-08 pvth0=6.904070074e-15 k1=7.583304170e-01 lk1=-3.083862960e-07 wk1=-5.385129682e-08 pk1=9.879262372e-14 k2=-1.206755324e-01 lk2=1.236130417e-07 wk2=1.969604640e-08 pk2=-3.907410513e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.928004152e-01 ldsub=6.722585984e-08 wdsub=7.267770858e-09 pdsub=-7.270612556e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.236767915e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.390485881e-07 wvoff=8.538058420e-08 pvoff=-6.383642673e-14 nfactor=-4.910563813e+00 lnfactor=6.178172271e-06 wnfactor=3.000995384e-06 pnfactor=-2.449217421e-12 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-1.561251128e-23 peta0=-2.081668171e-29 etab=-7.242729124e-01 letab=3.615889322e-07 wetab=2.398060949e-07 petab=-1.197734411e-13 u0=4.983145375e-02 lu0=-1.972601450e-08 wu0=-1.074422721e-08 pu0=7.048284447e-15 ua=8.724600159e-10 lua=-1.689913401e-15 wua=-7.205605234e-16 pua=5.894440746e-22 ub=7.327705034e-19 lub=9.264243670e-25 wub=2.635216704e-25 pub=-3.479364833e-31 uc=-1.528058854e-10 luc=1.825327169e-16 wuc=7.734960573e-17 puc=-7.310995813e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.369485432e+05 lvsat=2.137710017e-01 wvsat=1.639370697e-01 pvsat=-3.169741550e-8 a0=-5.904212609e-01 la0=7.970067687e-07 wa0=6.924353193e-07 pa0=-2.640021161e-13 ags=8.835138808e+00 lags=-4.116225816e-06 wags=-2.798990645e-06 pags=1.302865102e-12 a1=0.0 a2=0.42385546 b0=2.810164514e-06 lb0=-1.406181031e-12 wb0=-1.142424564e-12 pb0=5.716589699e-19 b1=-1.282966260e-08 lb1=6.419847697e-15 wb1=1.521613204e-14 pb1=-7.614015526e-21 keta=-6.338293872e-01 lketa=3.047138474e-07 wketa=2.223238947e-07 pketa=-1.074154643e-13 dwg=0.0 dwb=0.0 pclm=7.566914246e-01 lpclm=-4.332688117e-07 wpclm=2.296388946e-07 ppclm=6.144227363e-15 pdiblc1=6.652170123e-01 lpdiblc1=-1.089816360e-06 wpdiblc1=4.631194040e-09 ppdiblc1=3.312381736e-13 pdiblc2=6.005356984e-03 lpdiblc2=-5.101060662e-09 wpdiblc2=1.440829564e-09 ppdiblc2=1.929405464e-16 pdiblcb=4.894546198e-01 lpdiblcb=-4.076292767e-07 wpdiblcb=-1.704089772e-07 ppdiblcb=1.350239369e-13 drout=2.598793554e+00 ldrout=-8.000221209e-07 wdrout=-7.587483942e-07 pdrout=3.796709392e-13 pscbe1=1.796511879e+09 lpscbe1=-1.282076227e+03 wpscbe1=-3.300865878e+02 ppscbe1=4.246774937e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.258632522e-05 lalpha0=-8.884611950e-12 walpha0=-1.097297787e-11 palpha0=3.131986101e-18 alpha1=0.85 beta0=3.277913068e+01 lbeta0=-3.378489476e-06 wbeta0=-6.843622480e-06 pbeta0=1.696134939e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.181481947e-01 lkt1=1.411529985e-08 wkt1=-2.251639909e-08 pkt1=-7.940414242e-15 kt2=-6.558302836e-02 lkt2=3.626168475e-08 wkt2=2.072437873e-08 pkt2=-1.977921015e-14 at=-3.666661975e+05 lat=2.064694098e-01 wat=2.076118387e-01 pat=-1.115033245e-7 ute=-3.772240095e+00 lute=1.520720237e-06 wute=1.265041459e-06 pute=-7.575481371e-13 ua1=-5.819340951e-09 lua1=4.078960581e-15 wua1=3.256373200e-15 pua1=-1.953259957e-21 ub1=6.150856428e-18 lub1=-4.529205096e-24 wub1=-2.958203754e-24 pub1=1.969798128e-30 uc1=3.663556311e-10 luc1=-3.471601754e-16 wuc1=-1.250763042e-16 puc1=1.344800893e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.159 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='7.140932978e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.249969019e-08 wvth0=-3.761431814e-08 pvth0=9.418286734e-15 k1=-6.241904741e-01 lk1=3.834147152e-07 wk1=2.873836778e-07 pk1=-7.195828647e-14 k2=3.986372134e-01 lk2=-1.362463825e-07 wk2=-1.168735231e-07 pk2=2.926407833e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.954585123e-01 ldsub=6.589577199e-08 wdsub=-1.453554172e-08 pdsub=3.639568826e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236273e-03 lcdscd=-1.677929252e-09 wcdscd=-1.734723476e-24 pcdscd=4.336808690e-31 cit=0.0 voff='8.709368161e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.649725970e-08 wvoff=-8.445100331e-08 pvoff=2.114577117e-14 nfactor=1.294122777e+01 lnfactor=-2.754703571e-06 wnfactor=-3.790185361e-06 pnfactor=9.490283027e-13 eta0=9.800711343e-01 leta0=-2.452271850e-7 etab=4.074395393e-02 letab=-2.121862259e-08 wetab=8.934822982e-10 petab=-2.237199261e-16 u0=5.822572835e-04 lu0=4.917840169e-09 wu0=6.687879403e-09 pu0=-1.674584812e-15 ua=-3.900591379e-09 lua=6.984785594e-16 wua=9.155282949e-16 pua=-2.292400453e-22 ub=3.998140878e-18 lub=-7.075375803e-25 wub=-8.642904446e-25 pub=2.164105487e-31 uc=3.315753443e-10 luc=-5.984729108e-17 wuc=-1.376196463e-16 puc=3.445872085e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-2.533316142e+05 lvsat=1.218907430e-01 wvsat=2.013408750e-01 pvsat=-5.041394303e-8 a0=5.039151347e-01 la0=2.494106854e-07 wa0=3.299451431e-07 pa0=-8.261529432e-14 ags=-3.276249260e-02 lags=3.211921833e-07 wags=-3.908985055e-07 pags=9.787746768e-14 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.348334955e-02 lketa=-2.920344024e-08 wketa=1.533364699e-08 pketa=-3.839407205e-15 dwg=0.0 dwb=0.0 pclm=-4.574520557e-01 lpclm=1.742776586e-07 wpclm=4.842138539e-07 ppclm=-1.212427911e-13 pdiblc1=-3.385321472e+00 lpdiblc1=9.370366423e-07 wpdiblc1=1.334222326e-06 ppdiblc1=-3.340772623e-13 pdiblc2=-1.680339556e-02 lpdiblc2=6.312233832e-09 wpdiblc2=3.655674772e-09 ppdiblc2=-9.153480618e-16 pdiblcb=-5.473850359e-01 lpdiblcb=1.111959554e-07 wpdiblcb=1.990112736e-07 ppdiblcb=-4.983063181e-14 drout=1.497449274e+00 ldrout=-2.489193556e-07 wdrout=2.859143353e-13 pdrout=-7.159037629e-20 pscbe1=-2.325129067e+09 lpscbe1=7.803558074e+02 wpscbe1=1.038020544e+03 ppscbe1=-2.599110019e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.966353388e-05 lalpha0=-7.422073466e-12 walpha0=-9.435173069e-12 palpha0=2.362482420e-18 alpha1=0.85 beta0=3.775317354e+01 lbeta0=-5.867455757e-06 wbeta0=-6.913408631e-06 pbeta0=1.731055300e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.388387712e-01 lkt1=-2.557042189e-08 wkt1=-7.682967079e-08 pkt1=1.923745810e-14 kt2=4.270221610e-02 lkt2=-1.792327701e-08 wkt2=-3.763567022e-08 pkt2=9.423633103e-15 at=6.320637255e+04 lat=-8.634955368e-03 wat=-3.046491582e-02 pat=7.628140736e-9 ute=-1.463928423e-01 lute=-2.936210957e-07 wute=-4.981311058e-07 pute=1.247275457e-13 ua1=4.691943605e-09 lua1=-1.180791610e-15 wua1=-1.295200460e-15 pua1=3.243065383e-22 ub1=-6.514347683e-18 lub1=1.808349055e-24 wub1=1.958158372e-24 pub1=-4.903052330e-31 uc1=-8.027729087e-10 luc1=2.378612237e-16 wuc1=2.875721294e-16 puc1=-7.200547304e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.160 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='-1.170623630e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.392339810e-07 wvth0=2.288994019e-07 pvth0=-5.731435015e-14 k1=9.070734895e-01 lk1=8.724976297e-17 k2=-2.238942992e-01 lk2=1.962990551e-08 wk2=3.005524488e-08 pk2=-7.525562820e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.867948969e+00 ldsub=-3.528807861e-07 wdsub=-6.077575310e-07 pdsub=1.521770159e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999993e-03 lcdscd=1.357951945e-18 wcdscd=7.486702230e-19 pcdscd=-1.874605072e-25 cit=0.0 voff='-1.036177346e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.874483749e-08 wvoff=-9.807699097e-17 pvoff=2.455757819e-23 nfactor=-1.398124776e+01 lnfactor=3.986441999e-06 wnfactor=6.532145212e-06 pnfactor=-1.635590372e-12 eta0=2.482946376e-03 leta0=-4.479009417e-10 weta0=9.146675275e-16 peta0=-2.290245169e-22 etab=-4.399800002e-02 letab=3.767236523e-18 u0=-4.283222971e-02 lu0=1.578843698e-08 wu0=2.095300391e-08 pu0=-5.246443601e-15 ua=-1.910834825e-09 lua=2.002614262e-16 wua=2.954219006e-16 pua=-7.397098512e-23 ub=-1.524510109e-18 lub=6.752845231e-25 wub=6.700871844e-25 pub=-1.677838002e-31 uc=2.560381357e-10 luc=-4.093345388e-17 wuc=-5.321099410e-17 puc=1.332355402e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.091095223e+04 lvsat=4.070332254e-02 wvsat=5.726596730e-02 pvsat=-1.433888282e-8 a0=1.499999999e+00 la0=2.665325738e-16 ags=1.250000000e+00 lags=5.706635164e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.810340918e-01 lketa=1.246661964e-07 wketa=1.523111786e-07 pketa=-3.813734833e-14 dwg=0.0 dwb=0.0 pclm=4.071416362e-01 lpclm=-4.220882055e-08 wpclm=-6.823411541e-09 ppclm=1.708520839e-15 pdiblc1=3.569721503e-01 lpdiblc1=-4.562961120e-17 pdiblc2=8.406112093e-03 lpdiblc2=1.223434548e-18 pdiblcb=-1.032957700e-01 lpdiblcb=3.622435685e-18 drout=5.033266587e-01 ldrout=2.416733480e-16 pscbe1=7.914198799e+08 lpscbe1=2.387523651e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.843339998e-07 lalpha0=-4.074712889e-14 walpha0=-7.951279629e-14 palpha0=1.990928858e-20 alpha1=0.85 beta0=2.008012246e+01 lbeta0=-1.442282823e-06 wbeta0=-1.976283713e-06 pbeta0=4.948436553e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.740714101e-01 lkt1=-1.674848621e-08 wkt1=-3.922886275e-08 pkt1=9.822554174e-15 kt2=-2.887893901e-02 lkt2=1.448174913e-18 at=-1.210664066e+05 lat=3.750529007e-02 wat=3.681147971e-02 pat=-9.217263216e-9 ute=-1.014086739e+00 lute=-7.635835333e-08 wute=-1.351590028e-07 pute=3.384259787e-14 ua1=-2.384733751e-11 lua1=2.732435152e-25 ub1=7.077531678e-19 lub1=3.881553877e-34 uc1=1.471862500e-10 luc1=-5.620175274e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.161 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='1.455915859e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.255118363e-07 wvth0=-3.162445296e-07 pvth0=4.102470880e-14 k1=0.90707349 k2=-2.473606389e-02 lk2=-1.629644771e-08 wk2=-3.355345016e-08 pk2=3.948873287e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-7.388858263e-01 ldsub=1.173687496e-07 wdsub=4.513555915e-07 pdsub=-3.887745935e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000005e-03 lcdscd=-7.931294510e-19 wcdscd=-1.746897765e-18 pcdscd=2.627177989e-25 cit=0.0 voff='4.807727367e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.610925173e-08 wvoff=-8.466786455e-08 pvoff=1.527332076e-14 nfactor=4.850481829e+01 lnfactor=-7.285481942e-06 wnfactor=-1.879205364e-05 pnfactor=2.932667183e-12 eta0=-1.234617175e-02 leta0=2.227138684e-09 weta0=4.089571032e-09 peta0=-7.377218720e-16 etab=-0.043998 u0=1.028337804e-01 lu0=-1.048840024e-08 wu0=-3.627331928e-08 pu0=5.076670066e-15 ua=-1.565470016e-09 lua=1.379607228e-16 wua=2.148009587e-16 pua=-5.942769278e-23 ub=-4.262580240e-18 lub=1.169207732e-24 wub=8.122999829e-25 pub=-1.934377091e-31 uc=-5.073355809e-10 luc=9.677229424e-17 wuc=2.368801085e-16 puc=-3.900627006e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-8.013286645e+05 lvsat=1.980474992e-01 wvsat=2.931586747e-01 pvsat=-5.689180421e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.825838234e-02 lketa=2.675434341e-08 wketa=2.991628524e-08 pketa=-1.605841112e-14 dwg=0.0 dwb=0.0 pclm=-2.814011759e-02 lpclm=3.631209030e-08 wpclm=1.313961834e-07 ppclm=-2.322505011e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.002221418e-07 lalpha0=6.470153805e-14 walpha0=1.855298571e-13 palpha0=-2.790202072e-20 alpha1=0.85 beta0=3.235839949e+00 lbeta0=1.596274144e-06 wbeta0=4.611328657e-06 pbeta0=-6.935023278e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.970358441e-01 lkt1=2.347229101e-08 wkt1=9.153401338e-08 pkt1=-1.376589182e-14 kt2=-0.028878939 at=2.528974051e+05 lat=-2.995441588e-02 wat=-8.589345257e-02 pat=1.291760222e-8 ute=-1.895542474e+00 lute=8.264832816e-08 wute=1.045788211e-07 pute=-9.403947924e-15 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.162 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.163 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.647792282e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.431421449e-7 k1=5.566409778e-01 lk1=2.273392882e-7 k2=-2.306999056e-02 lk2=-1.959309392e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017412205e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.307349451e-7 nfactor=4.102012727e+00 lnfactor=-5.208356362e-6 eta0=0.08 etab=-0.07 u0=1.998563880e-02 lu0=2.504571366e-8 ua=-1.134300921e-09 lua=1.763046897e-15 wua=8.271806126e-31 ub=1.354178821e-18 lub=-8.817936668e-25 uc=6.336172452e-11 luc=-2.965002869e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.479005689e+00 la0=-2.328159296e-06 wa0=-8.881784197e-22 ags=3.213721844e-01 lags=4.701655027e-07 wags=-2.220446049e-22 a1=0.0 a2=0.42385546 b0=-1.166562766e-08 lb0=2.336724415e-13 wb0=1.809457590e-31 pb0=-3.670613968e-35 b1=1.188900229e-08 lb1=-2.822059756e-14 keta=-1.960740289e-03 lketa=-5.171820529e-8 dwg=0.0 dwb=0.0 pclm=-2.756450521e-02 lpclm=8.888074800e-07 ppclm=-2.220446049e-28 pdiblc1=0.39 pdiblc2=-1.582993035e-04 lpdiblc2=2.237297265e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.699568392e+07 lpscbe1=5.840027849e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.784862809e-01 lkt1=-1.578774688e-7 kt2=-2.846521888e-02 lkt2=-2.105465392e-8 at=1.883339850e+05 lat=-2.666849136e-1 ute=-1.123933750e+00 lute=1.706783447e-7 ua1=8.759880256e-10 lua1=4.900335287e-15 ub1=-2.475009312e-19 lub1=-6.439507266e-24 uc1=4.318848194e-11 luc1=-1.874060626e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.164 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.987799311e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=7.112322725e-8 k1=6.074244362e-01 lk1=-1.789482353e-7 k2=-5.399866830e-02 lk2=5.151057588e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.260430581e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.368925737e-8 nfactor=3.893743274e+00 lnfactor=-3.542119304e-6 eta0=0.08 etab=-0.07 u0=2.086568003e-02 lu0=1.800503969e-8 ua=-1.226154067e-09 lua=2.497907974e-15 ub=1.522777252e-18 lub=-2.230647031e-24 uc=3.260261592e-11 luc=-5.041539131e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.206001760e+00 la0=-1.440211147e-7 ags=4.067426001e-01 lags=-2.128312028e-7 a1=0.0 a2=0.42385546 b0=6.801093286e-08 lb0=-4.037711962e-13 wb0=-1.323488980e-29 pb0=1.058791184e-34 b1=6.982465203e-09 lb1=1.103361762e-14 keta=-1.930756365e-02 lketa=8.706316418e-08 wketa=-6.938893904e-24 dwg=0.0 dwb=0.0 pclm=-3.479201702e-01 lpclm=3.451778059e-06 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.070139653e-03 lpdiblc2=2.966805198e-8 pdiblcb=-0.025 drout=0.56 pscbe1=5.259308455e+08 lpscbe1=1.096383779e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.826384771e-01 lkt1=-1.246582759e-7 kt2=-1.849409519e-02 lkt2=-1.008275422e-7 at=1.700014663e+05 lat=-1.200175956e-1 ute=-8.049709096e-01 lute=-2.381149096e-6 ua1=2.398568951e-09 lua1=-7.280907441e-15 ub1=-1.692312545e-18 lub1=5.119550569e-24 uc1=-1.219150133e-11 luc1=2.556554572e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.165 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.083418339e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.287187748e-8 k1=5.214903467e-01 lk1=1.648217229e-7 k2=-2.253367664e-02 lk2=-7.436169359e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.116046597e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.930018581e-9 nfactor=2.923983519e+00 lnfactor=3.372988903e-7 eta0=0.08 etab=-0.07 u0=2.695731094e-02 lu0=-6.363865778e-9 ua=-5.110436127e-10 lua=-3.628134508e-16 ub=9.502970929e-19 lub=5.949744365e-26 uc=-5.459976453e-12 luc=1.018498607e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.198670600e+04 lvsat=2.720797692e-1 a0=8.399354850e-01 la0=1.320387115e-6 ags=4.387166488e-01 lags=-3.407398992e-7 a1=0.0 a2=0.42385546 b0=1.965027587e-08 lb0=-2.103096592e-13 pb0=5.293955920e-35 b1=-2.730237572e-09 lb1=4.988822639e-14 keta=-1.301593619e-02 lketa=6.189419433e-08 wketa=-3.469446952e-24 dwg=0.0 dwb=0.0 pclm=-7.677707209e-01 lpclm=5.131344424e-06 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=-7.243652152e-04 lpdiblc2=2.828481903e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.055883949e-01 lkt1=-3.284963096e-8 kt2=-5.695790970e-02 lkt2=5.304275524e-8 at=140000.0 ute=-1.615642111e+00 lute=8.618526807e-7 ua1=-3.363388199e-10 lua1=3.659792990e-15 ub1=6.699373247e-20 lub1=-1.918362431e-24 uc1=5.820842900e-11 luc1=-2.597179049e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.166 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.012513060e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.705570559e-8 k1=6.221540504e-01 lk1=-3.654504390e-8 k2=-6.385021927e-02 lk2=8.287546430e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.770949775e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.186573841e-8 nfactor=3.251393364e+00 lnfactor=-3.176488161e-7 eta0=1.574990403e-01 leta0=-1.550283827e-7 etab=-1.397147478e-01 letab=1.394567541e-7 u0=2.860688814e-02 lu0=-9.663665155e-9 ua=-1.713048856e-10 lua=-1.042423743e-15 ub=5.555140752e-19 lub=8.492178392e-25 uc=4.837013937e-11 luc=-5.831418567e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.199890520e+05 lvsat=5.603284828e-2 a0=1.5 ags=3.345158490e-01 lags=-1.322975571e-7 a1=0.0 a2=0.42385546 b0=1.483724021e-07 lb0=-4.678042421e-13 b1=2.787321384e-08 lb1=-1.133064239e-14 keta=1.805641432e-02 lketa=-2.626559775e-10 dwg=0.0 dwb=0.0 pclm=2.559697942e+00 lpclm=-1.524893942e-6 pdiblc1=1.905165224e-01 lpdiblc1=3.990449531e-7 pdiblc2=2.099520489e-02 lpdiblc2=-1.516281354e-8 pdiblcb=-0.025 drout=4.657394385e-01 ldrout=1.885579788e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.480538192e-01 lkt1=5.209782144e-8 kt2=-3.442621933e-02 lkt2=7.970564605e-9 at=1.500039100e+05 lat=-2.001173153e-2 ute=-1.650654028e+00 lute=9.318902044e-7 ua1=7.917739496e-10 lua1=1.403126358e-15 ub1=-4.209751012e-19 lub1=-9.422339682e-25 uc1=4.288729629e-11 luc1=4.676465496e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.167 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.241313638e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.416670170e-8 k1=5.957565380e-01 lk1=-1.013721011e-8 k2=-6.121433361e-02 lk2=5.650630147e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.147413854e-01 ldsub=4.527631070e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.591785940e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.366980730e-8 nfactor=4.149263696e+00 lnfactor=-1.215870216e-6 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-4.857225733e-23 peta0=-8.326672685e-29 etab=-0.0003125 u0=1.739526749e-02 lu0=1.552339234e-9 ua=-1.302869572e-09 lua=8.958338552e-17 ub=1.528326835e-18 lub=-1.239752905e-25 uc=8.070799787e-11 luc=-3.818192117e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.796777092e+04 lvsat=1.180783797e-1 a0=1.5 ags=3.851516517e-01 lags=-1.829531584e-7 a1=0.0 a2=0.42385546 b0=-6.387476527e-07 lb0=3.196235767e-13 b1=3.310693975e-08 lb1=-1.656641469e-14 keta=3.735329723e-02 lketa=-1.956708397e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=1.449957661e+00 lpclm=-4.147197528e-07 wpclm=-8.881784197e-22 pdiblc1=6.791983131e-01 lpdiblc1=-8.982791209e-8 pdiblc2=1.035513619e-02 lpdiblc2=-4.518584568e-9 pdiblcb=-0.025 drout=3.081770429e-01 ldrout=3.461819813e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.404457400e-07 lalpha0=5.706687843e-13 walpha0=-5.293955920e-29 palpha0=-2.646977960e-35 alpha1=0.85 beta0=1.211863932e+01 lbeta0=1.742041552e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.861238714e-01 lkt1=-9.856340949e-9 kt2=-3.017355137e-03 lkt2=-2.345058046e-8 at=2.601016600e+05 lat=-1.301525297e-1 ute=4.684522305e-02 lute=-7.662727686e-7 ua1=4.011457076e-09 lua1=-1.817815664e-15 ub1=-2.779785683e-18 lub1=1.417498909e-24 uc1=-1.124233100e-11 luc1=5.882725747e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.168 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='7.381111596e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.495029008e-07 wvth0=1.744740323e-07 pvth0=-8.730523552e-14 k1=2.434038474e-01 lk1=1.661769051e-07 wk1=-4.504498996e-16 pk1=2.254010312e-22 k2=-2.347538467e-03 lk2=-2.380578434e-08 wk2=1.594946806e-08 pk2=-7.980970273e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.812004566e+00 ldsub=-7.539798094e-07 wdsub=-5.500034896e-07 pdsub=2.752167962e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236286e-03 lcdscd=-1.677929258e-09 wcdscd=-4.089013850e-18 pcdscd=2.046106340e-24 cit=0.0 voff='-4.600177942e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.435342532e-07 wvoff=9.677529615e-08 pvoff=-4.842548722e-14 nfactor=-1.332830712e+01 lnfactor=7.529748924e-06 wnfactor=4.911387916e-06 pnfactor=-2.457614311e-12 eta0=9.730901924e-01 leta0=-2.417339358e-07 weta0=2.312413398e-09 peta0=-1.157110853e-15 etab=4.344132419e-02 letab=-2.189401984e-08 wetab=-1.944930675e-17 petab=9.732272930e-24 u0=1.998912111e-02 lu0=2.543982305e-10 wu0=2.595110163e-10 pu0=-1.298569770e-16 ua=-1.495965753e-09 lua=1.862069768e-16 wua=1.190152934e-16 pua=-5.955418170e-23 ub=4.019133765e-18 lub=-1.370352661e-24 wub=-8.712441703e-25 pub=4.359627416e-31 uc=-9.496309798e-11 luc=4.972231416e-17 wuc=3.667800435e-18 puc=-1.835334327e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.142158131e+05 lvsat=-1.014583439e-02 wvsat=1.334533009e-02 pvsat=-6.677883069e-9 a0=1.500000005e+00 la0=-2.285734269e-15 wa0=-1.376042391e-15 pa0=6.885589876e-22 ags=-1.212861952e+00 lags=6.166784668e-07 wags=-2.946227984e-16 pags=1.474265363e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.283382739e-01 lketa=-1.151342474e-07 wketa=-4.921048785e-08 pketa=2.462448522e-14 dwg=0.0 dwb=0.0 pclm=4.268819652e-01 lpclm=9.721811755e-08 wpclm=1.912852841e-07 ppclm=-9.571743460e-14 pdiblc1=6.426167888e-01 lpdiblc1=-7.152284655e-08 wpdiblc1=2.355755591e-16 ppdiblc1=-1.178798170e-22 pdiblc2=-5.767129694e-03 lpdiblc2=3.548852181e-09 wpdiblc2=-6.316313791e-18 ppdiblc2=3.160626275e-24 pdiblcb=5.341822465e-02 lpdiblcb=-3.923977385e-08 wpdiblcb=-1.870215094e-17 ppdiblcb=9.358375186e-24 drout=1.497450141e+00 ldrout=-2.489195736e-07 wdrout=-1.247705050e-15 pdrout=6.243403572e-22 pscbe1=8.085935397e+08 lpscbe1=-4.300129932e+00 wpscbe1=-1.232633591e-07 ppscbe1=6.167960167e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.481017758e-06 lalpha0=-4.408533568e-13 walpha0=-9.994006402e-14 palpha0=5.000910857e-20 alpha1=0.85 beta0=1.768657030e+01 lbeta0=-1.044101000e-06 wbeta0=-2.665068398e-07 pbeta0=1.333576241e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.696409066e-01 lkt1=-6.814336819e-08 wkt1=-6.662670987e-08 pkt1=3.333940598e-14 kt2=-7.091764556e-02 lkt2=1.052611377e-08 wkt2=-7.476519404e-18 pkt2=3.741187915e-24 at=1.220911654e+05 lat=-6.109332034e-02 wat=-4.997003237e-02 pat=2.500455447e-8 ute=-1.247936989e+00 lute=-1.183754027e-07 wute=-1.332534196e-07 pute=6.667881188e-14 ua1=7.818100525e-10 lua1=-2.017293603e-16 wua1=-1.410693669e-24 pua1=7.058983572e-31 ub1=-6.027834062e-19 lub1=3.281465622e-25 wub1=-2.003958322e-33 pub1=1.002762714e-39 uc1=6.539033548e-11 luc1=2.048096086e-17 wuc1=2.901594492e-26 puc1=-1.451934620e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.169 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='2.560494590e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.731402609e-07 wvth0=-6.231215441e-07 pvth0=1.124055185e-13 k1=9.070734847e-01 lk1=9.633591702e-16 wk1=1.608750466e-15 pk1=-2.902040830e-22 k2=3.880677982e-02 lk2=-3.411045525e-08 wk2=-5.696238594e-08 pk2=1.027550176e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-5.896935037e+00 ldsub=1.176269287e-06 wdsub=1.964298177e-06 pdsub=-3.543417125e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999952e-03 lcdscd=8.745002986e-18 wcdscd=1.460362387e-17 pcdscd=-2.634362346e-24 cit=0.0 voff='9.398068842e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.069692479e-07 wvoff=-3.456260577e-07 pvoff=6.234783017e-14 nfactor=5.869316050e+01 lnfactor=-1.050377838e-05 wnfactor=-1.754067113e-05 pnfactor=3.164179206e-12 eta0=2.741523461e-02 leta0=-4.945461092e-09 weta0=-8.258619278e-09 peta0=1.489780590e-15 etab=-4.399800023e-02 letab=4.159544931e-17 wetab=6.946188069e-17 petab=-1.253029625e-23 u0=2.322167941e-02 lu0=-5.550052752e-10 wu0=-9.268250584e-10 pu0=1.671908991e-16 ua=2.642411619e-10 lua=-2.545329929e-16 wua=-4.250546195e-16 pua=7.667602786e-23 ub=-8.895251555e-18 lub=1.863293194e-24 wub=3.111586323e-24 pub=-5.613021683e-31 uc=1.349432660e-10 luc=-7.844170233e-18 wuc=-1.309928727e-17 puc=2.362993529e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.876819549e+05 lvsat=-2.854109511e-02 wvsat=-4.766189318e-02 pvsat=8.597776572e-9 a0=1.499999984e+00 la0=2.942883270e-15 wa0=4.914433305e-15 pa0=-8.865197465e-22 ags=1.249999997e+00 lags=6.300968636e-16 wags=1.052224974e-15 pags=-1.898121660e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.517997666e-01 lketa=1.052443967e-07 wketa=1.757517423e-07 pketa=-3.170403255e-14 dwg=0.0 dwb=0.0 pclm=2.448967001e+00 lpclm=-4.090937766e-07 wpclm=-6.831617289e-07 ppclm=1.232362274e-13 pdiblc1=3.569721528e-01 lpdiblc1=-5.038152118e-16 wpdiblc1=-8.413403307e-16 ppdiblc1=1.517702630e-22 pdiblc2=8.406112025e-03 lpdiblc2=1.350843049e-17 wpdiblc2=2.255826081e-17 ppdiblc2=-4.069303922e-24 pdiblcb=-1.032957702e-01 lpdiblcb=3.999744980e-17 wpdiblcb=6.679345965e-17 ppdiblcb=-1.204894517e-23 drout=5.033266452e-01 ldrout=2.668414822e-15 wdrout=4.456090608e-15 pdrout=-8.038387733e-22 pscbe1=7.914198785e+08 lpscbe1=2.636175156e-07 wpscbe1=4.402236938e-07 ppscbe1=-7.941246033e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.133257357e-06 lalpha0=2.137376036e-13 walpha0=3.569288001e-13 palpha0=-6.438674317e-20 alpha1=0.85 beta0=1.124038035e+01 lbeta0=5.699669481e-07 wbeta0=9.518101423e-07 pbeta0=-1.716979834e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.010865651e+00 lkt1=1.424917368e-07 wkt1=2.379525352e-07 pkt1=-4.292449578e-14 kt2=-2.887893909e-02 lkt2=1.598970956e-17 wkt2=2.670186294e-17 pkt2=-4.816778920e-24 at=-5.487081960e+05 lat=1.068688026e-01 wat=1.784644013e-01 pat=-3.219337182e-8 ute=-2.858853021e+00 lute=2.849834734e-07 wute=4.759050700e-07 pute=-8.584899148e-14 ua1=-2.384735272e-11 lua1=3.016991073e-24 wua1=5.038191623e-24 pua1=-9.088444257e-31 ub1=7.077531462e-19 lub1=4.285781150e-33 wub1=7.156994489e-33 pub1=-1.291057346e-39 uc1=1.471862503e-10 luc1=-6.205508955e-26 wuc1=-1.036283600e-25 puc1=1.869366146e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.170 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='-6.434254564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.048180802e-07 wvth0=3.791454863e-07 pvth0=-6.839443341e-14 k1=0.90707349 k2=-1.051417275e-01 lk2=-8.143440074e-09 wk2=-6.919717345e-09 pk2=1.248254732e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.427842290e+00 ldsub=-5.058366201e-07 wdsub=-9.288397632e-07 pdsub=1.675543337e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='4.807716122e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.610923142e-08 wvoff=-8.466782730e-08 pvoff=1.527331403e-14 nfactor=2.491112224e+00 lnfactor=-3.654346851e-07 wnfactor=-3.550381611e-06 pnfactor=6.404568892e-13 eta0=0.0 etab=-0.043998 u0=3.623981224e-02 lu0=-2.903359274e-09 wu0=-1.421460009e-08 pu0=2.564185925e-15 ua=-3.646487008e-09 lua=4.509271723e-16 wua=9.041211891e-16 pua=-1.630953254e-22 ub=-8.982807731e-18 lub=1.879087540e-24 wub=2.375837577e-24 pub=-4.285797164e-31 uc=-1.191640290e-10 luc=3.799449883e-17 wuc=1.083013873e-16 puc=-1.953659556e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-9.854663233e+05 lvsat=2.191624960e-01 wvsat=3.541528011e-01 pvsat=-6.388597795e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.111168377e+00 lketa=1.881103596e-07 wketa=3.853091375e-07 pketa=-6.950630063e-14 dwg=0.0 dwb=0.0 pclm=1.992526528e-02 lpclm=2.908349112e-08 wpclm=1.154749098e-07 ppclm=-2.083063446e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.598815119e-07 lalpha0=-1.953301020e-14 walpha0=2.698696521e-21 palpha0=-4.868205662e-28 alpha1=0.85 beta0=1.715716828e+01 lbeta0=-4.973683427e-07 wbeta0=1.866987986e-14 pbeta0=-3.367880197e-21 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.207000705e-01 lkt1=-1.808612243e-08 wkt1=-9.297602688e-16 pkt1=1.677203931e-22 kt2=-0.028878939 at=-6.409845432e+03 lat=9.043060798e-03 wat=-2.986065811e-10 pat=5.386595149e-17 ute=-9.684077382e-01 lute=-5.603584160e-08 wute=-2.025271429e-07 pute=3.653407383e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.171 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.481936+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.032866346 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.8416 eta0=0.08 etab=-0.07 u0=0.0212379 ua=-1.0461503e-9 ub=1.31009e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=1.7766e-11 b1=1.0478e-8 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.172 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.647792282e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.431421449e-7 k1=5.566409778e-01 lk1=2.273392882e-7 k2=-2.306999056e-02 lk2=-1.959309392e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017412205e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.307349451e-07 wvoff=-5.551115123e-23 nfactor=4.102012727e+00 lnfactor=-5.208356362e-6 eta0=0.08 etab=-0.07 u0=1.998563880e-02 lu0=2.504571366e-8 ua=-1.134300921e-09 lua=1.763046897e-15 ub=1.354178821e-18 lub=-8.817936668e-25 uc=6.336172452e-11 luc=-2.965002869e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.479005689e+00 la0=-2.328159296e-06 wa0=-8.881784197e-22 ags=3.213721844e-01 lags=4.701655027e-7 a1=0.0 a2=0.42385546 b0=-1.166562766e-08 lb0=2.336724415e-13 wb0=-3.218249571e-30 pb0=7.237830360e-36 b1=1.188900229e-08 lb1=-2.822059756e-14 keta=-1.960740289e-03 lketa=-5.171820529e-8 dwg=0.0 dwb=0.0 pclm=-2.756450521e-02 lpclm=8.888074800e-7 pdiblc1=0.39 pdiblc2=-1.582993035e-04 lpdiblc2=2.237297265e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.699568392e+07 lpscbe1=5.840027849e+03 ppscbe1=9.536743164e-19 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.784862809e-01 lkt1=-1.578774688e-7 kt2=-2.846521888e-02 lkt2=-2.105465392e-8 at=1.883339850e+05 lat=-2.666849136e-1 ute=-1.123933750e+00 lute=1.706783447e-7 ua1=8.759880256e-10 lua1=4.900335287e-15 ub1=-2.475009312e-19 lub1=-6.439507266e-24 uc1=4.318848194e-11 luc1=-1.874060626e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.173 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='4.987799311e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=7.112322725e-8 k1=6.074244362e-01 lk1=-1.789482353e-7 k2=-5.399866830e-02 lk2=5.151057588e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.260430581e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.368925737e-8 nfactor=3.893743274e+00 lnfactor=-3.542119304e-6 eta0=0.08 etab=-0.07 u0=2.086568003e-02 lu0=1.800503969e-8 ua=-1.226154067e-09 lua=2.497907974e-15 ub=1.522777252e-18 lub=-2.230647031e-24 uc=3.260261592e-11 luc=-5.041539131e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.206001759e+00 la0=-1.440211147e-7 ags=4.067426002e-01 lags=-2.128312028e-7 a1=0.0 a2=0.42385546 b0=6.801093286e-08 lb0=-4.037711962e-13 pb0=-5.293955920e-35 b1=6.982465203e-09 lb1=1.103361762e-14 keta=-1.930756365e-02 lketa=8.706316418e-08 wketa=-6.938893904e-24 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=-3.479201702e-01 lpclm=3.451778059e-06 wpclm=5.551115123e-23 ppclm=2.220446049e-28 pdiblc1=0.39 pdiblc2=-1.070139653e-03 lpdiblc2=2.966805198e-08 ppdiblc2=6.938893904e-30 pdiblcb=-0.025 drout=0.56 pscbe1=5.259308455e+08 lpscbe1=1.096383779e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.826384771e-01 lkt1=-1.246582759e-7 kt2=-1.849409519e-02 lkt2=-1.008275422e-7 at=1.700014663e+05 lat=-1.200175956e-1 ute=-8.049709096e-01 lute=-2.381149096e-6 ua1=2.398568951e-09 lua1=-7.280907441e-15 ub1=-1.692312545e-18 lub1=5.119550569e-24 uc1=-1.219150133e-11 luc1=2.556554572e-16 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.174 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.083418339e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.287187748e-8 k1=5.214903467e-01 lk1=1.648217229e-7 k2=-2.253367664e-02 lk2=-7.436169359e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.116046597e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.930018581e-9 nfactor=2.923983519e+00 lnfactor=3.372988903e-7 eta0=0.08 etab=-0.07 u0=2.695731094e-02 lu0=-6.363865778e-9 ua=-5.110436127e-10 lua=-3.628134508e-16 ub=9.502970929e-19 lub=5.949744365e-26 uc=-5.459976452e-12 luc=1.018498607e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.198670600e+04 lvsat=2.720797692e-1 a0=8.399354850e-01 la0=1.320387115e-6 ags=4.387166488e-01 lags=-3.407398992e-7 a1=0.0 a2=0.42385546 b0=1.965027587e-08 lb0=-2.103096592e-13 b1=-2.730237572e-09 lb1=4.988822639e-14 keta=-1.301593619e-02 lketa=6.189419433e-8 dwg=0.0 dwb=0.0 pclm=-7.677707209e-01 lpclm=5.131344424e-6 pdiblc1=0.39 pdiblc2=-7.243652152e-04 lpdiblc2=2.828481903e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.055883949e-01 lkt1=-3.284963096e-8 kt2=-5.695790970e-02 lkt2=5.304275524e-8 at=140000.0 ute=-1.615642111e+00 lute=8.618526807e-7 ua1=-3.363388199e-10 lua1=3.659792990e-15 pua1=8.271806126e-37 ub1=6.699373247e-20 lub1=-1.918362431e-24 uc1=5.820842900e-11 luc1=-2.597179049e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.175 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.012513060e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.705570559e-8 k1=6.221540504e-01 lk1=-3.654504390e-8 k2=-6.385021927e-02 lk2=8.287546430e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.601173000e-01 ldsub=-6.003519459e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.770949775e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.186573841e-8 nfactor=3.251393364e+00 lnfactor=-3.176488161e-7 eta0=1.574990403e-01 leta0=-1.550283827e-7 etab=-1.397147478e-01 letab=1.394567541e-7 u0=2.860688814e-02 lu0=-9.663665155e-9 ua=-1.713048856e-10 lua=-1.042423743e-15 ub=5.555140752e-19 lub=8.492178392e-25 uc=4.837013937e-11 luc=-5.831418567e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.199890520e+05 lvsat=5.603284828e-2 a0=1.5 ags=3.345158490e-01 lags=-1.322975571e-7 a1=0.0 a2=0.42385546 b0=1.483724021e-07 lb0=-4.678042421e-13 pb0=1.058791184e-34 b1=2.787321384e-08 lb1=-1.133064239e-14 keta=1.805641432e-02 lketa=-2.626559775e-10 dwg=0.0 dwb=0.0 pclm=2.559697942e+00 lpclm=-1.524893942e-6 pdiblc1=1.905165224e-01 lpdiblc1=3.990449531e-7 pdiblc2=2.099520489e-02 lpdiblc2=-1.516281354e-8 pdiblcb=-0.025 drout=4.657394385e-01 ldrout=1.885579788e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.480538192e-01 lkt1=5.209782144e-8 kt2=-3.442621933e-02 lkt2=7.970564605e-9 at=1.500039100e+05 lat=-2.001173153e-2 ute=-1.650654028e+00 lute=9.318902044e-7 ua1=7.917739496e-10 lua1=1.403126358e-15 ub1=-4.209751012e-19 lub1=-9.422339682e-25 uc1=4.288729629e-11 luc1=4.676465496e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.176 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='5.241313638e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.416670170e-8 k1=5.957565380e-01 lk1=-1.013721011e-8 k2=-6.121433361e-02 lk2=5.650630147e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.147413854e-01 ldsub=4.527631070e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.591785940e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.366980730e-8 nfactor=4.149263696e+00 lnfactor=-1.215870216e-6 eta0=-4.853187006e-01 leta0=4.880406999e-07 weta0=-6.938893904e-24 peta0=-9.194034423e-29 etab=-0.0003125 u0=1.739526749e-02 lu0=1.552339234e-9 ua=-1.302869572e-09 lua=8.958338552e-17 ub=1.528326835e-18 lub=-1.239752905e-25 uc=8.070799787e-11 luc=-3.818192117e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.796777092e+04 lvsat=1.180783797e-1 a0=1.5 ags=3.851516517e-01 lags=-1.829531584e-07 wags=2.220446049e-22 a1=0.0 a2=0.42385546 b0=-6.387476527e-07 lb0=3.196235767e-13 b1=3.310693975e-08 lb1=-1.656641469e-14 keta=3.735329723e-02 lketa=-1.956708397e-8 dwg=0.0 dwb=0.0 pclm=1.449957661e+00 lpclm=-4.147197528e-7 pdiblc1=6.791983131e-01 lpdiblc1=-8.982791209e-8 pdiblc2=1.035513619e-02 lpdiblc2=-4.518584568e-9 pdiblcb=-0.025 drout=3.081770429e-01 ldrout=3.461819813e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.404457400e-07 lalpha0=5.706687843e-13 walpha0=5.293955920e-29 palpha0=1.323488980e-35 alpha1=0.85 beta0=1.211863932e+01 lbeta0=1.742041552e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-2.861238714e-01 lkt1=-9.856340949e-9 kt2=-3.017355137e-03 lkt2=-2.345058046e-8 at=2.601016600e+05 lat=-1.301525297e-1 ute=4.684522305e-02 lute=-7.662727686e-7 ua1=4.011457076e-09 lua1=-1.817815664e-15 ub1=-2.779785683e-18 lub1=1.417498909e-24 uc1=-1.124233100e-11 luc1=5.882725747e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.177 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='6.529934091e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.031470602e-8 k1=2.434038459e-01 lk1=1.661769059e-7 k2=5.059815988e-02 lk2=-5.029933529e-08 pk2=-1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.378164456e-02 ldsub=1.596271782e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.753236272e-03 lcdscd=-1.677929251e-9 cit=0.0 voff='-1.387634666e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.721852107e-8 nfactor=2.975488218e+00 lnfactor=-6.285235302e-7 eta0=9.807663600e-01 leta0=-2.455750696e-7 etab=4.344132412e-02 letab=-2.189401981e-08 wetab=-2.385244779e-24 petab=1.355252716e-30 u0=2.085059134e-02 lu0=-1.766737215e-10 ua=-1.100883748e-09 lua=-1.148850293e-17 ub=1.126960129e-18 lub=7.686499680e-26 uc=-8.278750349e-11 luc=4.362975626e-17 puc=8.077935669e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.585168405e+05 lvsat=-3.231366978e-2 a0=1.5 ags=-1.212861953e+00 lags=6.166784673e-07 wags=-1.387778781e-23 pags=-4.857225733e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.497961921e-02 lketa=-3.339104685e-08 wketa=-3.469446952e-24 pketa=-1.734723476e-30 dwg=0.0 dwb=0.0 pclm=1.061870725e+00 lpclm=-2.205245432e-7 pdiblc1=6.426167896e-01 lpdiblc1=-7.152284695e-8 pdiblc2=-5.767129715e-03 lpdiblc2=3.548852191e-09 ppdiblc2=-2.168404345e-31 pdiblcb=5.341822458e-02 lpdiblcb=-3.923977382e-8 drout=1.497450137e+00 ldrout=-2.489195716e-7 pscbe1=8.085935393e+08 lpscbe1=-4.300129728e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.149257698e-06 lalpha0=-2.748436086e-13 alpha1=0.85 beta0=1.680187680e+01 lbeta0=-6.014083338e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-3.908142817e-01 lkt1=4.252979816e-8 kt2=-7.091764558e-02 lkt2=1.052611378e-8 at=-4.378886584e+04 lat=2.191155437e-2 ute=-1.690283739e+00 lute=1.029709298e-7 ua1=7.818100478e-10 lua1=-2.017293580e-16 ub1=-6.027834128e-19 lub1=3.281465655e-25 wub1=9.629649722e-41 pub1=3.611118646e-47 uc1=6.539033558e-11 luc1=2.048096081e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.178 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='0.4919864+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.90707349 k2=-0.150285 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.62373 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=0.46532 eta0=0.0 etab=-0.043998 u0=0.020145 ua=-1.146766e-9 ub=1.43394e-18 uc=9.1459e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=229464.0 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.068376 dwg=0.0 dwb=0.0 pclm=0.18115 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.16e-8 alpha1=0.85 beta0=14.4 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=43720.487 ute=-1.2790432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.179 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.299402e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0365*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=4.4379e-8 lint=-1.955e-10 vth0='-5.761948103e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.926902767e-07 wvth0=3.588927920e-07 pvth0=-6.474102964e-14 k1=0.90707349 k2=-2.127292966e-01 lk2=1.126438910e-08 wk2=2.549017715e-08 pk2=-4.598198546e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.348307880e+00 ldsub=-4.914893283e-07 wdsub=-9.048806583e-07 pdsub=1.632323268e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='4.807717192e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.610923335e-08 wvoff=-8.466783052e-08 pvoff=1.527331462e-14 nfactor=2.491112037e+00 lnfactor=-3.654346514e-07 wnfactor=-3.550381555e-06 pnfactor=6.404568790e-13 eta0=0.0 etab=-0.043998 u0=-1.079238621e-01 lu0=2.310247010e-08 wu0=2.921355350e-08 pu0=-5.269862129e-15 ua=-3.646487209e-09 lua=4.509272086e-16 wua=9.041212498e-16 pua=-1.630953364e-22 ub=-8.982836031e-18 lub=1.879092645e-24 wub=2.375846103e-24 pub=-4.285812543e-31 uc=-1.098904349e-10 luc=3.632162591e-17 wuc=1.055077913e-16 puc=-1.903265597e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.545278688e+05 lvsat=1.351780364e-02 wvsat=1.073867070e-02 pvsat=-1.937159546e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.111168044e+00 lketa=1.881102996e-07 wketa=3.853090373e-07 pketa=-6.950628255e-14 dwg=0.0 dwb=0.0 pclm=1.992536747e-02 lpclm=2.908347269e-08 wpclm=1.154748791e-07 ppclm=-2.083062891e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.598815202e-07 lalpha0=-1.953301170e-14 walpha0=1.949577618e-22 palpha0=-3.516859621e-29 alpha1=0.85 beta0=1.715716834e+01 lbeta0=-4.973683538e-07 wbeta0=3.410605132e-17 pbeta0=-6.153300092e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=-6.13e-10 dwc=2.252e-8 xpart=0.0 cgso=2.4892e-10 cgdo=2.4892e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.00154845795 mjs=0.44 pbsws=0.2 cjsws=4.24559793e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.75331171e-10 mjswgs=0.8 tnom=30.0 kt1=-1.207000734e-01 lkt1=-1.808612191e-08 wkt1=-7.255618328e-17 pkt1=1.308853026e-23 kt2=-0.028878939 at=-6.409846347e+03 lat=9.043060963e-03 wat=-2.302019857e-11 pat=4.152621841e-18 ute=-9.857496776e-01 lute=-5.290751180e-08 wute=-1.973030224e-07 pute=3.559168951e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.ends sky130_fd_pr__nfet_01v8