* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_pfet_01v8_b__toxe_mult=0.948
.param sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult=0.8
.param sky130_fd_pr__rf_pfet_01v8_b__overlap_mult=0.95436
.param sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult=0.90161
.param sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult=0.90587
.param sky130_fd_pr__rf_pfet_01v8_b__lint_diff=1.7325e-8
.param sky130_fd_pr__rf_pfet_01v8_b__wint_diff=-3.2175e-8
.param sky130_fd_pr__rf_pfet_01v8_b__rshg_diff=-7.0
.param sky130_fd_pr__rf_pfet_01v8_b__dlc_diff=1.7325e-8
.param sky130_fd_pr__rf_pfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__xgw_diff=-6.4250e-8
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult=0.85
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult=0.77
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult=0.77
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2=0.85
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2=0.80
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2=0.80
.param sky130_fd_pr__rf_pfet_01v8__aw_rd_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rs_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_0=0.0036576
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_0=-0.00034614
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_0=-0.092407
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_0=-19636.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_1=-0.0076806
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_1=-0.00019683
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_1=-0.079373
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_1=-15546.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_2=-0.033345
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_2=-3.0791e-5
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_2=-0.030098
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_2=-6434.1
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_3=-0.0012925
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_3=-0.00028011
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_3=-0.12131
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_3=-18686.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_4=0.00024736
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_4=-0.00041476
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_4=-0.071611
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_4=-11333.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_5=-0.016582
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_5=-0.00016695
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_5=-0.025831
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_5=-1107.2
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_6=-0.0014721
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_6=-0.00053506
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_6=-0.13112
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_6=-16484.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_7=-0.00025473
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_7=-17993.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_7=0.00033491
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_7=-0.077674
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_8=-0.035077
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_8=-0.00020922
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_8=-5719.7
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_8=-0.019564
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_0=0.0065905
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_0=-0.00050702
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_0=-0.081008
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_0=-20196.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_1=-0.0063812
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_1=-0.00027314
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_1=-0.065695
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_1=-12293.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_2=-7.2735e-5
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_2=-0.022778
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_2=272.66
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_2=-0.034415
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_3=0.00078898
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_3=-0.0003818
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_3=-0.11908
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_3=-16139.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_4=-0.00058216
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_4=-0.058416
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_4=-11485.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_4=0.0039762
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_5=-0.01803
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_5=-0.00025609
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_5=-7303.4
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_5=-0.016473
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_6=-0.12568
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_6=-0.00035343
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_6=-16543.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_6=0.00030278
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_7=0.0028314
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_7=-0.073523
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_7=-0.000511
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_7=-15224.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_8=-0.018202
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_8=-0.022497
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_8=-0.00030626
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_8=4136.5
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_8=0.0
.include "sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"