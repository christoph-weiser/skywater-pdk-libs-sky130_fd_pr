* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult=1.0365
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult=1.2
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult=9.6320e-1
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult=1.1229e+0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult=1.0009e+0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff=-1.21275e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff=2.252e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff=7.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff=-1.1228e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff=4.504e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42=1.1125
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42=1.245
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42=1.245
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult=1.1125
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult=1.245
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult=1.245
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_0=0.035472
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_0=-0.0035791
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_0=11669.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_0=-0.023208
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_1=-0.015447
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_1=0.031659
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_1=-0.0022517
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_1=16627.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_2=-0.00027242
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_2=0.006014
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_2=-0.0024036
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_2=7476.5
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_3=-0.025698
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_3=0.022412
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_3=-0.0067063
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_3=14950.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_4=-0.018667
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_4=0.0074967
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_4=-0.0031604
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_4=14641.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_5=-0.0050153
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_5=0.005408
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_5=-0.0036655
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_5=14592.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_6=-0.031185
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_6=0.019026
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_6=-0.0097006
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_6=9042.7
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_7=-0.018406
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_7=0.005177
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_7=-0.0054184
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_7=13962.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_8=-0.0045172
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_8=0.0026993
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_8=-0.0049523
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_8=16409.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_0=-0.022384
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_0=0.032174
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_0=-0.0088162
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_0=18475.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_1=-0.015672
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_1=0.024627
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_1=-0.0052084
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_1=17204.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_2=-0.0053553
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_2=0.00058529
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_2=-0.0047533
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_2=14144.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_3=-0.026679
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_3=0.025797
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_3=-0.0070348
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_3=14175.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_4=-0.007826
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_4=18436.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_4=-0.019062
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_4=0.0093971
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_5=-0.0078718
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_5=-0.0066522
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_5=26781.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_5=-0.0060231
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_6=-0.03107
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_6=0.017691
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_6=-0.0077169
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_6=12148.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_7=-0.019933
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_7=0.0024544
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_7=-0.0097882
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_7=13883.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_8=-0.0057624
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_8=-0.0093065
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_8=39684.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_8=-0.014919
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_8=0.0
.include "sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"