* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_g5v0d16v0__toxe_mult=0.9635
.param sky130_fd_pr__pfet_g5v0d16v0__rshp_mult=1.0
.param sky130_fd_pr__pfet_g5v0d16v0__soverlap_mult=0.40
.param sky130_fd_pr__pfet_g5v0d16v0__doverlap_mult=0.40
.param sky130_fd_pr__pfet_g5v0d16v0__ajunction_mult=9.5405e-1
.param sky130_fd_pr__pfet_g5v0d16v0__pjunction_mult=9.6374e-1
.param sky130_fd_pr__pfet_g5v0d16v0__wint_diff=-2.252e-8
.param sky130_fd_pr__pfet_g5v0d16v0__lint_diff=1.21275e-8
.param sky130_fd_pr__pfet_g5v0d16v0__dlc_diff=1.21275e-8
.param sky130_fd_pr__pfet_g5v0d16v0__dwc_diff=-2.252e-88
.param sky130_fd_pr__pfet_g5v0d16v0__cf_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cjswgs_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigc_diff=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdiff_mult=0.6024
.param sky130_fd_pr__pfet_g5v0d16v0__aigbinv_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ua_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbacc_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nigbacc_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__dsub_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bigsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__a0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__lpe0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigc_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__keta_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ub_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__k2_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ags_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vth0_diff_0=0.041
.param sky130_fd_pr__pfet_g5v0d16v0__u0_diff_0=3.6814e-3
.param sky130_fd_pr__pfet_g5v0d16v0__nigbinv_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__voff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__jtssws_diff_0=-4.02e-12
.param sky130_fd_pr__pfet_g5v0d16v0__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__voff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbinv_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ua_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigbacc_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nigbacc_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__dsub_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bigsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__aigsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__a0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__lpe0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__keta_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ub_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__k2_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__ags_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__vth0_diff_1=1.2588e-2
.param sky130_fd_pr__pfet_g5v0d16v0__u0_diff_1=4.0038e-3
.param sky130_fd_pr__pfet_g5v0d16v0__nigbinv_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__b1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d16v0__jtssws_diff_1=-4.02e-12