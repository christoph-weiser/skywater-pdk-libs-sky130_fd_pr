* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__special_nfet_pass_lvt__toxe_mult=1.0
.param sky130_fd_pr__special_nfet_pass_lvt__overlap_mult=9.2429e-1
.param sky130_fd_pr__special_nfet_pass_lvt__ajunction_mult=1.0004e+0
.param sky130_fd_pr__special_nfet_pass_lvt__pjunction_mult=8.9176e-1
.param sky130_fd_pr__special_nfet_pass_lvt__rshn_mult=1.0
.param sky130_fd_pr__special_nfet_pass_lvt__lint_diff=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__wint_diff=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__dlc_diff=-1.3619e-9
.param sky130_fd_pr__special_nfet_pass_lvt__dwc_diff=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__u0_diff_0=-6.9731e-3
.param sky130_fd_pr__special_nfet_pass_lvt__vsat_diff_0=8.1112e+3
.param sky130_fd_pr__special_nfet_pass_lvt__vth0_diff_0=2.4767e-2
.param sky130_fd_pr__special_nfet_pass_lvt__nfactor_diff_0=4.0502e-1
.param sky130_fd_pr__special_nfet_pass_lvt__voff_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__k2_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__ua_diff_0=0.0
.param sky130_fd_pr__special_nfet_pass_lvt__ub_diff_0=0.0
.include "sky130_fd_pr__special_nfet_pass_lvt.pm3.spice"