* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param tol_nfom=-0.0483u
.param tol_pfom=-0.042u
.param tol_nw=-0.0483u
.param tol_poly=-0.0287u
.param tol_li=-0.014u
.param tol_m1=-0.0175u
.param tol_m2=-0.0175u
.param tol_m3=-0.0455u
.param tol_m4=-0.0455u
.param tol_m5=-0.119u
.param tol_rdl=-0.7u
.param rcn=296.1
.param rcp=789
.param rdn=128.4
.param rdp=218.7
.param rdn_hv=122.4
.param rdp_hv=212.7
.param rp1=53.52
.param rnw=2022
.param rl1=14.02
.param rm1=0.139
.param rm2=0.139
.param rm3=0.0533
.param rm4=0.0533
.param rm5=0.03361
.param rrdl=0.00617
.param rcp1=213.88
.param rcl1=18.61
.param rcvia=11.85
.param rcvia2=6.623
.param rcvia3=6.623
.param rcvia4=0.7377
.param rcrdlcon=0.00713
.param rspwres=4120
.param crpf_precision=1.39e-04
.param crpfsw_precision_1_1=5.59e-11
.param crpfsw_precision_2_1=5.95e-11
.param crpfsw_precision_4_1=6.41e-11
.param crpfsw_precision_8_2=6.96e-11
.param crpfsw_precision_16_2=7.61e-11
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/slow_70p.spice"