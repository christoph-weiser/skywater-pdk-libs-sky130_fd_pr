* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_hvt__toxe_mult=1.0
.param sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_hvt__overlap_mult=0.98867
.param sky130_fd_pr__pfet_01v8_hvt__lint_diff=0.0
.param sky130_fd_pr__pfet_01v8_hvt__wint_diff=0.0
.param sky130_fd_pr__pfet_01v8_hvt__dlc_diff=0.0
.param sky130_fd_pr__pfet_01v8_hvt__dwc_diff=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=0.64787
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=-0.11577
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=-0.00842
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=9.171e-20
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.00036389
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=-7112.2
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=0.026419
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=-1.6478246e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=3.7374e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=-0.16912
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=-0.1709
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=0.6412
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=-0.12187
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=-2.2902e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=-0.016292
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.0010687
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=-7333.7
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=0.011671
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=-6.7051481e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=3.4586e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=0.20802
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=0.0096114
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=-0.014652
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=-0.038521
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=3.8706e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=-0.0057008
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0015318
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=-0.011385
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=-4.933e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=-4.6376e-11
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=-1.9658e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=0.28726
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=0.00017109
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=-0.00015832
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=-0.026013
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=3.2924e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=-0.0085614
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.001453
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.003849
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=-1.1139e-10
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=-1.7119e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=-7.2896e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=0.21396
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=-0.026141
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.032133
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=-0.040491
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=3.5687e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=-0.0098132
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.001225
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=-0.000998
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=1.2597e-8
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=-3.4893e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=0.26111
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=0.037081
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=-0.040342
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=-0.042255
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=3.6307e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=-0.010815
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.0015534
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=-0.0012997
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=-5.3637136e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=3.469e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=-0.15276
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=0.96493
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=-0.17885
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=-2.4224e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=-0.025463
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0012069
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=-1169.8
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=0.00010707
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=-0.00071726
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=5.0661e-19
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=58018.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=-0.018827
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=-2.2466963e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=-4.5014e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.046706
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=0.68647
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=-0.14245
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=-0.0029197
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=-0.0052868
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=-0.00016947
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=-7.4084e-20
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=5.5373
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=-0.0067962
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=-1.5741e-11
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=1.6004e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=0.94739
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=-0.13932
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=-0.042856
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=-0.009604
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0014206
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=2.5647e-19
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=43211.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.00081692
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=-1.7966e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=5.7833e-11
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=0.11217
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=2.4575e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=-0.038563
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=0.026757
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=-0.036831
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=-1.8971e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=0.14974
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.00080614
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.0030218
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=-0.013242
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=-5.8082e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=-3.411e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=6.2077e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=-0.047257
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=0.00061775
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=-0.0010307
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=-1.0557e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=0.21755
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.0001177
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=0.0070281
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=-0.014467
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=-0.003503
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=-1.1408e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=1.847e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=0.00017941
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=-0.031808
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=0.022826
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=-3.5419e-12
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=1.1994
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.00013703
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=0.0096373
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=1.2343
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=-1.4672e-5
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=0.020459
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=-0.005387
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=-1.1232e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=-2.0802e-21
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=-0.0079777
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=-0.038083
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=0.024895
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=-1.0198e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=-10064.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=0.54598
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.00039043
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=0.024758
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=-0.01124
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=3.7828e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=7.0659e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=-0.20026
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=-0.095719
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=-1.3101263e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=36284.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=0.90538
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.00054452
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=-0.01158
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=-0.013393
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=-1.4565e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=2.0802e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.15162
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=-0.16446
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=-3.2055002e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=-6011.3
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=0.78817
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.00036165
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=-0.014737
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0064619
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=5.6362e-12
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=1.7598e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=-0.10862
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=-8.3152e-11
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=-5.9285e-11
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=1.2823
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=-6.2466e-6
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=28075.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.0080941
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=-0.0031058
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=-1.1089e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=4.2583e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=-0.021129
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=0.046321
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=-0.066616
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=-1.4484e-12
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=0.066563
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0013661
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=-0.0009615
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=-0.011723
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=-9.6778e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=4.4102e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=-0.040201
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=-0.044717
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.09561
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=-0.054159
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=-2.4008e-11
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=0.16473
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0012133
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=-0.0061071
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=-0.0077911
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=-2.0191e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=5.2225e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=-0.037085
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.059684
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=-0.0352
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=8.8703e-8
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=0.2151
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.00191
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=-0.0068057
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=-0.0071071
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=-1.9209e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=6.3617e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=6.067e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.1
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=-0.04099
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=0.002408
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=-0.0022284
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=4.0865e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=-0.36321
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=-0.0010792
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.011949
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=-0.0044603
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=-6.1271e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=4.0977e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=2.7114e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=-0.13858
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=-0.087652
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=-1.0e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=-12916.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=0.45894
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=0.00034876
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=0.0088449
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=-0.011624
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=-0.0073835
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=1.6227e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=7.6056e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.16014
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=-0.13917
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=-1.0e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=20012.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=0.78898
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.0010815
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=0.0063494
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=0.92326
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.00035054
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=-0.017067
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=-0.0045308
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=-5.212e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=2.6633e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=-0.12196
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=-6.4121e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=12736.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=44084.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=-0.33053
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=-1.5871e-5
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.0066354
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=-0.0099005
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=-1.5878e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=2.6336e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=-0.03415
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=-8.318e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=-0.00032957
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0018413
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=-0.0067644
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=-0.0095046
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=-1.4936e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=5.6221e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=-0.044741
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.093361
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=-0.0643
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=-6.012e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=0.089097
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.0018157
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=-0.0032836
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=-0.007636
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=-1.7667e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=5.8807e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=-0.030487
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.084638
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=-0.049385
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=-9.4896e-11
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=-1.2144e-10
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=1.2166
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0014352
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.0091372
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=-0.0053636
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=-1.3672e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=2.9847e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=-0.0059034
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=0.016143
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=-0.0093132
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=0.0032384
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=-0.0026603
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=-6.6748e-12
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=1.2187
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0017419
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.0035912
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=-0.0088595
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=-1.4852e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=3.3671e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=-0.0078252
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=-0.079774
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=-6596.7
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=0.52228
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.0012291
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=0.0026861
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=-0.029749
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=3.1813e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=-1.8716e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=-0.21153
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.16741
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=-0.15643
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=-1.0e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=25963.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=0.9368
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=0.00014681
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=-0.022563
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=-0.011281
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=-1.4225e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=3.0833e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=1.6451e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.15
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=-0.032636
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=-4.5646e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=3307.1
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=0.12366
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.00016422
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=-0.0052903
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=-0.0028117
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=-1.7243e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=-2.4885e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=2.5424e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=-0.01298
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=-7.0533e-11
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=31234.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=1.2891
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0010899
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=-0.0053108
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=-0.010171
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=-0.0031312
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=-2.371e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=3.4376e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=-0.054193
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=-1.087e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=-6.4382e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=2.1543e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=1.387
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0014966
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=-0.012619
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=0.22953
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.0021307
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=-0.044111
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=-0.009361
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=-1.4456e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=5.2005e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=-0.055437
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=-1.8059e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=-8.9873e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=3.3859e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=1.2381
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=-0.00032659
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=0.015101
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=0.0069385
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=-9.0008e-12
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=-2.4281e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=-0.01182
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=-1.9465e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=3.6662e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=8.0158e-8
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=1.8873e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=0.22912
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0020212
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=-0.021515
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=-0.0055742
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=-1.3629e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=5.3159e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=-0.050147
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=-1.4529e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=-5.1926e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=-1.9645e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=7.79e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=1.2423
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.00064866
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=-0.014047
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=-0.0019647
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=-2.527e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=9.7792e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=-0.015728
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=-7.1716e-10
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=-4.1396435e-9
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=0.75251
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.00046506
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=2353.7
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.040283
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=-0.0064094
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=7.7102e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=8.1554e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=-0.33699
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=-0.18153
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=-2.9262738e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=35823.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=0.70173
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=-0.00097972
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.026116
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=-0.0075535
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=-4.8538e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=4.9561e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=-0.067496
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=-0.19665
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=-0.040166
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=-9.9273e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=23057.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=1.4109
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.00077483
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.029596
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=-0.010991
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=-2.5485e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=2.1997e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=-0.06677
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=-1.2236e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=-9.9363e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=3.1242e-8
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=0.29746
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0021119
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=-0.019842
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=-0.010603
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=1.1179e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=2.6904e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=3.8482e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=-0.042159
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=-8.099e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=-4.0065e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=2.1896e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=0.27193
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.0013084
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=-0.0037886
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=-0.0028399
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=-5.5028e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=-8.7318e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=4.68e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=-0.046546
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=-3.6266e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=-7.0024e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=1.8226e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=0.29301
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0018674
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=-0.011215
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=-0.0048261
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=0.00053147
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=-4.9698e-12
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=-3.4539e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=-0.017283
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=-5.0381e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=3.1378e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=2.9495e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=0.088947
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=-5.6365e-5
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.020368
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=0.43295
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.00071
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=-0.011557
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=-0.02751
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=1.5449e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=-2.8376e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=-0.10752
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=-0.11006
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=-1.0698583e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=8644.1
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=-13180.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=1.3992
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.00092803
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.017853
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=-0.0026549
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=1.1727e-12
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=2.7682e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=-0.03499
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=-8.9529e-10
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=5438.5
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=0.80855
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=-3.1814e-5
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=0.018002
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=-0.0084157
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=-8.6721e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=1.5947e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=-0.19977
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=-0.17477
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=-1.035337e-9
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=-6586.5
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=0.60686
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.00018862
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=0.049411
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=-0.01019
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=-7.9353e-12
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=7.604e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=-0.30131
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=-0.11721
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=-1.03534e-9
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=16.90778869
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=0.00248037
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=-0.19976997
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=-0.08250904
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=-1.31013e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=189.96735041
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=3.13009e-6
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.25855998
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=-0.00076997
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=-0.20025994
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=-0.054395
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=-0.09801202
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=-5.36378e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=-109.76124038
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=-1.3001e-6
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=-0.16616984
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=0.00030941
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=-0.15275999
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=-0.17090007
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=-0.089626
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=-6.70515e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=93.10299601
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=1.30003e-6
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=0.03262997
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=-0.00024997
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=-0.30130994
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=-0.06820702
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=-439.92974224
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=-4.20007e-6
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=-0.80763995
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=0.00125002
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.15162
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=-0.10678
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=-3.2055e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=3360.00200157
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=1.19797e-5
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=0.77924005
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=-0.0026698
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=-0.020934
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=-0.11116
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=81981.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=-0.00017582
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.020045
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=-0.00017618
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.77573
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=0.0019559
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=-0.014348
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=78372.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=36202.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=-0.00020189
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=1.0141
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=0.0061561
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=-0.015801
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=25602.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=-0.00016346
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=0.9613
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=0.0020874
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=-0.014445
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=25454.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=-0.0001819
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=0.77033
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=0.0013599
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=-0.013785
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=36053.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=-0.00021998
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=0.62741
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=0.0010395
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=-0.013308
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=37969.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=-0.00022145
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=0.68037
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=0.0025101
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=-0.011949
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=27669.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=-0.00015603
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=1.0832
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=0.0048176
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=-0.0098916
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=-0.24495
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=58607.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=-0.00011722
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=-0.0052133
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=-0.0068897
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=-0.44556
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=51004.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=-0.00031453
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.0014366
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=-0.0073046
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=52818.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=-0.0002412
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=0.71035
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=0.0022707
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=-0.012563
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=-0.01279
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=64603.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=-0.00029595
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=0.77624
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=0.0054188
.include "sky130_fd_pr__pfet_01v8_hvt.pm3.spice"