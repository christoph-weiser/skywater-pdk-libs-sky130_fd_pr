* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_lvt__toxe_mult=0.948
.param sky130_fd_pr__pfet_01v8_lvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_lvt__overlap_mult=0.1
.param sky130_fd_pr__pfet_01v8_lvt__ajunction_mult=9.0161e-1
.param sky130_fd_pr__pfet_01v8_lvt__pjunction_mult=9.0587e-1
.param sky130_fd_pr__pfet_01v8_lvt__lint_diff=1.7325e-8
.param sky130_fd_pr__pfet_01v8_lvt__wint_diff=-3.2175e-8
.param sky130_fd_pr__pfet_01v8_lvt__dlc_diff=3.417e-8
.param sky130_fd_pr__pfet_01v8_lvt__dwc_diff=-3.2175e-8
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_0=-0.00018181
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_0=-0.027802
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_0=0.10552
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_0=0.15965
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_0=0.076345
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_1=0.047725
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_1=-0.00011454
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_1=-0.01536
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_1=0.11088
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_1=0.13638
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_2=0.15683
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_2=0.051573
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_2=-0.00019763
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_2=-0.1008
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_2=0.11906
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_3=0.14152
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_3=0.053319
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_3=-0.00011326
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_3=-0.057942
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_3=0.11315
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_4=0.11569
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_4=4.3243e-8
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_4=0.069072
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_4=-0.00044707
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_4=-10072.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_4=2.0324e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_5=0.19325
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_5=4.3678e-7
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_5=0.062426
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_5=-0.00036688
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_5=-30803.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_5=4.8211e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_6=0.11742
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_6=0.08882
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_6=0.075834
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_6=0.045314
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_6=-0.00041292
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_7=1.0e-11
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_7=0.065344
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_7=0.076201
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_7=0.10547
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_7=0.072684
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_7=-0.00030377
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_8=0.0722
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_8=0.13399
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_8=0.088953
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_8=0.054843
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_8=-0.00046671
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_9=0.076126
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_9=0.12574
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_9=0.091349
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_9=0.057052
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_9=-0.0004448
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_10=-0.00043232
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_10=0.12887
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_10=0.046843
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_10=0.022448
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_10=0.10081
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_11=-0.00062778
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_11=-9231.3
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_11=0.094172
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_11=0.061969
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_12=0.03622
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_12=0.095072
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_12=-0.00055341
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_12=-20408.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_12=0.10158
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_12=-2.1123e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_13=0.053063
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_13=-0.090817
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_13=0.11048
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_13=-0.00036912
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_13=0.12098
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_14=0.048684
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_14=-0.10432
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_14=0.14664
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_14=-0.00026795
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_14=0.087931
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_15=0.062225
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_15=-0.067675
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_15=0.12282
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_15=-0.00043606
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_15=0.1536
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_16=0.062053
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_16=-0.016589
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_16=0.10606
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_16=-0.0003498
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_16=0.13219
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_17=0.051446
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_17=0.0033532
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_17=0.10371
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_17=-0.00035493
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_17=0.12997
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_18=0.052676
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_18=-0.00040195
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_18=-19653.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_18=0.071101
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_19=4.4057e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_19=0.035594
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_19=0.11429
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_19=-0.00039861
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_19=-24564.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_19=0.084123
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_20=0.039246
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_20=0.015874
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_20=0.14374
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_20=-0.00031632
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_20=0.08913
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_21=-0.0003466
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_21=0.083708
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_21=9.0e-12
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_21=0.063216
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_21=-0.029212
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_21=0.12512
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_22=0.08947
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_22=0.099093
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_22=-0.00026634
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_22=0.086469
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__uc_diff_22=1.3e-11
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_22=0.069371
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_23=0.053051
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_23=-0.055065
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_23=0.11871
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_23=-0.00029927
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_23=0.12288
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_24=0.050637
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_24=-0.033177
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_24=0.11867
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_24=-0.00026959
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_24=0.1185
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_25=0.049261
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_25=-0.00038249
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_25=-7742.9
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_25=0.040595
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_26=0.037948
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_26=0.09606
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_26=-0.00036152
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_26=-19903.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_26=0.073767
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_26=-7.8239e-8
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_27=1.8807e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_27=4.5094e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_27=0.07298
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_27=7.1187e-5
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_27=0.083832
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_27=-8.0e-3
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_28=1.6301e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_28=2.5833e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_28=0.026264
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_28=-0.00027633
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_28=0.088571
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_29=1.15e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_29=2.1875e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_29=0.042705
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_29=-0.00026294
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_29=0.13557
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_30=6.4792e-8
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_30=2.2441e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_30=0.045828
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_30=-0.00025477
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_30=0.10383
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_31=1.4677e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_31=1.8441e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_31=0.049127
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_31=-0.00032319
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_31=0.14753
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_32=-0.00027067
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_32=-21638.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_32=0.17994
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_32=0.07014
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_33=-0.00039943
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_33=-21782.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_33=0.13762
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_33=1.4751e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_33=2.0999e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_33=0.050551
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_34=0.074715
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_34=-0.00026303
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_34=0.15243
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_34=3.2237e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_34=5.0e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_35=0.065048
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_35=-0.00019647
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_35=0.12947
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_35=1.865e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_35=2.1007e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_36=0.069908
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_36=-0.00021967
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_36=0.12845
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_36=2.2594e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_36=2.0328e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_37=2.1218e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_37=0.051554
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_37=-0.00025681
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_37=0.10817
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_37=1.74e-7
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_38=0.05612
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_38=-0.00019302
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_38=-10913.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_38=0.052629
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_lvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b0_diff_39=2.3872e-7
.param sky130_fd_pr__pfet_01v8_lvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__b1_diff_39=3.8314e-7
.param sky130_fd_pr__pfet_01v8_lvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ub_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__k2_diff_39=0.046113
.param sky130_fd_pr__pfet_01v8_lvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__u0_diff_39=-0.00011531
.param sky130_fd_pr__pfet_01v8_lvt__vsat_diff_39=-27603.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_diff_39=0.077259
.param sky130_fd_pr__pfet_01v8_lvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_lvt__ua_diff_39=0.0
.include "sky130_fd_pr__pfet_01v8_lvt.pm3.spice"