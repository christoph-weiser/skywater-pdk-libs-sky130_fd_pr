* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8__toxe_mult=1.0365
.param sky130_fd_pr__pfet_01v8__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8__overlap_mult=1.1043
.param sky130_fd_pr__pfet_01v8__ajunction_mult=1.0625
.param sky130_fd_pr__pfet_01v8__pjunction_mult=1.0675
.param sky130_fd_pr__pfet_01v8__lint_diff=-1.21275e-8
.param sky130_fd_pr__pfet_01v8__wint_diff=2.252e-8
.param sky130_fd_pr__pfet_01v8__dlc_diff=-1.21275e-8
.param sky130_fd_pr__pfet_01v8__dwc_diff=2.252e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_0=-0.065212
.param sky130_fd_pr__pfet_01v8__vsat_diff_0=-6125.4
.param sky130_fd_pr__pfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_0=3.8528e-11
.param sky130_fd_pr__pfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_0=-0.023864
.param sky130_fd_pr__pfet_01v8__vth0_diff_0=0.051716
.param sky130_fd_pr__pfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_0=0.00025511
.param sky130_fd_pr__pfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_0=0.010183
.param sky130_fd_pr__pfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_0=1.6231e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_1=1.7969e-19
.param sky130_fd_pr__pfet_01v8__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_1=-0.16643
.param sky130_fd_pr__pfet_01v8__vsat_diff_1=-11757.0
.param sky130_fd_pr__pfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_1=2.6071e-11
.param sky130_fd_pr__pfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_1=-0.02798
.param sky130_fd_pr__pfet_01v8__vth0_diff_1=0.0095625
.param sky130_fd_pr__pfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_1=0.00048935
.param sky130_fd_pr__pfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_1=-0.012504
.param sky130_fd_pr__pfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_2=-0.038666
.param sky130_fd_pr__pfet_01v8__ags_diff_2=-0.085151
.param sky130_fd_pr__pfet_01v8__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_2=1.5678e-19
.param sky130_fd_pr__pfet_01v8__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_2=0.15084
.param sky130_fd_pr__pfet_01v8__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_2=0.091966
.param sky130_fd_pr__pfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_2=1.3913e-11
.param sky130_fd_pr__pfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_2=-0.011035
.param sky130_fd_pr__pfet_01v8__vth0_diff_2=-0.019558
.param sky130_fd_pr__pfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_2=0.00071619
.param sky130_fd_pr__pfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_3=-0.042662
.param sky130_fd_pr__pfet_01v8__ags_diff_3=0.017403
.param sky130_fd_pr__pfet_01v8__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_3=1.3946e-19
.param sky130_fd_pr__pfet_01v8__nfactor_diff_3=0.05285
.param sky130_fd_pr__pfet_01v8__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_3=-0.020048
.param sky130_fd_pr__pfet_01v8__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_3=-5.8266e-12
.param sky130_fd_pr__pfet_01v8__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_3=-0.012691
.param sky130_fd_pr__pfet_01v8__vth0_diff_3=-0.011216
.param sky130_fd_pr__pfet_01v8__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_3=0.00032572
.param sky130_fd_pr__pfet_01v8__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_4=0.00032453
.param sky130_fd_pr__pfet_01v8__vth0_diff_4=-0.021893
.param sky130_fd_pr__pfet_01v8__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_4=-0.038612
.param sky130_fd_pr__pfet_01v8__ags_diff_4=-0.016854
.param sky130_fd_pr__pfet_01v8__ub_diff_4=1.1269e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_4=0.040373
.param sky130_fd_pr__pfet_01v8__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_4=0.019253
.param sky130_fd_pr__pfet_01v8__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_4=7.4109e-13
.param sky130_fd_pr__pfet_01v8__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_4=-0.013076
.param sky130_fd_pr__pfet_01v8__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_5=-0.0094402
.param sky130_fd_pr__pfet_01v8__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_5=0.00019069
.param sky130_fd_pr__pfet_01v8__vth0_diff_5=-0.017541
.param sky130_fd_pr__pfet_01v8__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_5=-0.027577
.param sky130_fd_pr__pfet_01v8__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_5=0.0095471
.param sky130_fd_pr__pfet_01v8__ub_diff_5=7.2283e-20
.param sky130_fd_pr__pfet_01v8__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_5=0.016774
.param sky130_fd_pr__pfet_01v8__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_5=-0.0088631
.param sky130_fd_pr__pfet_01v8__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_5=-2.6578e-12
.param sky130_fd_pr__pfet_01v8__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_6=-0.033184
.param sky130_fd_pr__pfet_01v8__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_6=0.0003127
.param sky130_fd_pr__pfet_01v8__vth0_diff_6=-0.022738
.param sky130_fd_pr__pfet_01v8__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_6=0.0083827
.param sky130_fd_pr__pfet_01v8__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_6=1.6239e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_6=-0.096185
.param sky130_fd_pr__pfet_01v8__vsat_diff_6=3962.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_6=6.7557e-12
.param sky130_fd_pr__pfet_01v8__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_7=-5.7329e-11
.param sky130_fd_pr__pfet_01v8__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_7=-0.024181
.param sky130_fd_pr__pfet_01v8__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_7=-0.0001174
.param sky130_fd_pr__pfet_01v8__vth0_diff_7=-0.026431
.param sky130_fd_pr__pfet_01v8__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_7=-0.0015874
.param sky130_fd_pr__pfet_01v8__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_7=1.6007e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_7=-0.04787
.param sky130_fd_pr__pfet_01v8__vsat_diff_7=39789.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_8=8.1126e-11
.param sky130_fd_pr__pfet_01v8__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_8=-0.012783
.param sky130_fd_pr__pfet_01v8__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_8=-0.00090468
.param sky130_fd_pr__pfet_01v8__vth0_diff_8=0.0052319
.param sky130_fd_pr__pfet_01v8__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_8=0.015428
.param sky130_fd_pr__pfet_01v8__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_8=6.0112e-21
.param sky130_fd_pr__pfet_01v8__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_8=0.34648
.param sky130_fd_pr__pfet_01v8__vsat_diff_8=-35394.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_9=4.2884e-12
.param sky130_fd_pr__pfet_01v8__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_9=-0.011672
.param sky130_fd_pr__pfet_01v8__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_9=0.00036241
.param sky130_fd_pr__pfet_01v8__vth0_diff_9=0.0034908
.param sky130_fd_pr__pfet_01v8__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_9=-0.020849
.param sky130_fd_pr__pfet_01v8__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_9=1.159e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_9=0.048495
.param sky130_fd_pr__pfet_01v8__vsat_diff_9=-7053.8
.param sky130_fd_pr__pfet_01v8__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_10=37317.0
.param sky130_fd_pr__pfet_01v8__u0_diff_10=0.0015136
.param sky130_fd_pr__pfet_01v8__vth0_diff_10=-0.030253
.param sky130_fd_pr__pfet_01v8__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_10=-2.2543e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_10=0.2527
.param sky130_fd_pr__pfet_01v8__ub_diff_10=7.3478e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_10=-0.030257
.param sky130_fd_pr__pfet_01v8__voff_diff_10=-0.067326
.param sky130_fd_pr__pfet_01v8__a0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_11=-0.025163
.param sky130_fd_pr__pfet_01v8__a0_diff_11=0.030284
.param sky130_fd_pr__pfet_01v8__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_11=18141.0
.param sky130_fd_pr__pfet_01v8__u0_diff_11=0.0012435
.param sky130_fd_pr__pfet_01v8__vth0_diff_11=-0.027313
.param sky130_fd_pr__pfet_01v8__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_11=-2.0027e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_11=0.025446
.param sky130_fd_pr__pfet_01v8__ub_diff_11=3.4977e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_11=-0.02144
.param sky130_fd_pr__pfet_01v8__k2_diff_11=-0.015874
.param sky130_fd_pr__pfet_01v8__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_12=-0.018089
.param sky130_fd_pr__pfet_01v8__k2_diff_12=-0.012179
.param sky130_fd_pr__pfet_01v8__voff_diff_12=-0.024506
.param sky130_fd_pr__pfet_01v8__a0_diff_12=0.023887
.param sky130_fd_pr__pfet_01v8__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_12=0.0017386
.param sky130_fd_pr__pfet_01v8__vth0_diff_12=-0.021564
.param sky130_fd_pr__pfet_01v8__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_12=1.2332e-14
.param sky130_fd_pr__pfet_01v8__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_12=0.03969
.param sky130_fd_pr__pfet_01v8__ub_diff_12=4.3106e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_13=0.037538
.param sky130_fd_pr__pfet_01v8__ub_diff_13=4.1385e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_13=-0.0094728
.param sky130_fd_pr__pfet_01v8__k2_diff_13=-0.010252
.param sky130_fd_pr__pfet_01v8__voff_diff_13=-0.026089
.param sky130_fd_pr__pfet_01v8__a0_diff_13=0.012275
.param sky130_fd_pr__pfet_01v8__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_13=0.00168
.param sky130_fd_pr__pfet_01v8__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_13=-0.011631
.param sky130_fd_pr__pfet_01v8__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_13=-1.3656e-12
.param sky130_fd_pr__pfet_01v8__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_14=-1.0297e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_14=0.01182
.param sky130_fd_pr__pfet_01v8__ub_diff_14=3.6128e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_14=-0.02937
.param sky130_fd_pr__pfet_01v8__k2_diff_14=-0.0093488
.param sky130_fd_pr__pfet_01v8__voff_diff_14=-0.014191
.param sky130_fd_pr__pfet_01v8__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_14=0.039605
.param sky130_fd_pr__pfet_01v8__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_14=0.0014987
.param sky130_fd_pr__pfet_01v8__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_14=-0.007906
.param sky130_fd_pr__pfet_01v8__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_15=2.5233e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_15=-0.06052
.param sky130_fd_pr__pfet_01v8__ub_diff_15=2.3792e-19
.param sky130_fd_pr__pfet_01v8__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_15=-0.022612
.param sky130_fd_pr__pfet_01v8__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_15=-0.015348
.param sky130_fd_pr__pfet_01v8__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_15=0.00066818
.param sky130_fd_pr__pfet_01v8__vsat_diff_15=-15532.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_15=0.013505
.param sky130_fd_pr__pfet_01v8__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_16=3.0542e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_16=0.1063
.param sky130_fd_pr__pfet_01v8__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_16=2.3719e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_16=-0.021795
.param sky130_fd_pr__pfet_01v8__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_16=-0.024188
.param sky130_fd_pr__pfet_01v8__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_16=0.00071992
.param sky130_fd_pr__pfet_01v8__vsat_diff_16=-4787.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_16=0.018662
.param sky130_fd_pr__pfet_01v8__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_17=0.18027
.param sky130_fd_pr__pfet_01v8__ua_diff_17=2.3608e-11
.param sky130_fd_pr__pfet_01v8__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_17=3.1564e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_17=-0.013142
.param sky130_fd_pr__pfet_01v8__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_17=-0.01755
.param sky130_fd_pr__pfet_01v8__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_17=0.00049162
.param sky130_fd_pr__pfet_01v8__vsat_diff_17=-928.84
.param sky130_fd_pr__pfet_01v8__vth0_diff_17=-0.019812
.param sky130_fd_pr__pfet_01v8__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_18=0.27444
.param sky130_fd_pr__pfet_01v8__ua_diff_18=1.6549e-11
.param sky130_fd_pr__pfet_01v8__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_18=1.7799e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_18=-0.017655
.param sky130_fd_pr__pfet_01v8__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_18=-0.014193
.param sky130_fd_pr__pfet_01v8__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_18=0.00068138
.param sky130_fd_pr__pfet_01v8__vsat_diff_18=-20698.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_18=-0.011736
.param sky130_fd_pr__pfet_01v8__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_19=0.30807
.param sky130_fd_pr__pfet_01v8__ua_diff_19=2.0599e-11
.param sky130_fd_pr__pfet_01v8__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_19=-0.13971
.param sky130_fd_pr__pfet_01v8__ub_diff_19=2.9397e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_19=-0.0095155
.param sky130_fd_pr__pfet_01v8__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_19=-0.0074856
.param sky130_fd_pr__pfet_01v8__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_19=0.17095
.param sky130_fd_pr__pfet_01v8__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_19=0.0012038
.param sky130_fd_pr__pfet_01v8__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_19=-0.0039105
.param sky130_fd_pr__pfet_01v8__u0_diff_20=0.001381
.param sky130_fd_pr__pfet_01v8__vth0_diff_20=-0.011454
.param sky130_fd_pr__pfet_01v8__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_20=-1.4037e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_20=0.039603
.param sky130_fd_pr__pfet_01v8__ub_diff_20=3.5386e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_20=-0.011381
.param sky130_fd_pr__pfet_01v8__k2_diff_20=-0.014136
.param sky130_fd_pr__pfet_01v8__voff_diff_20=-0.021962
.param sky130_fd_pr__pfet_01v8__a0_diff_20=0.01444
.param sky130_fd_pr__pfet_01v8__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_21=0.0017077
.param sky130_fd_pr__pfet_01v8__vth0_diff_21=-0.0076811
.param sky130_fd_pr__pfet_01v8__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_21=-7.7891e-13
.param sky130_fd_pr__pfet_01v8__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_21=0.063402
.param sky130_fd_pr__pfet_01v8__ub_diff_21=3.7954e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_21=-0.044124
.param sky130_fd_pr__pfet_01v8__k2_diff_21=-0.013544
.param sky130_fd_pr__pfet_01v8__voff_diff_21=-0.023819
.param sky130_fd_pr__pfet_01v8__a0_diff_21=0.054291
.param sky130_fd_pr__pfet_01v8__voff_diff_22=-0.020991
.param sky130_fd_pr__pfet_01v8__a0_diff_22=0.052104
.param sky130_fd_pr__pfet_01v8__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_22=0.0018204
.param sky130_fd_pr__pfet_01v8__vth0_diff_22=-0.010234
.param sky130_fd_pr__pfet_01v8__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_22=-1.9323e-13
.param sky130_fd_pr__pfet_01v8__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_22=0.041898
.param sky130_fd_pr__pfet_01v8__ub_diff_22=4.0224e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_22=-0.042064
.param sky130_fd_pr__pfet_01v8__k2_diff_22=-0.013937
.param sky130_fd_pr__pfet_01v8__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_23=-0.017848
.param sky130_fd_pr__pfet_01v8__voff_diff_23=-0.024633
.param sky130_fd_pr__pfet_01v8__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_23=-11554.0
.param sky130_fd_pr__pfet_01v8__u0_diff_23=0.00072192
.param sky130_fd_pr__pfet_01v8__vth0_diff_23=0.025799
.param sky130_fd_pr__pfet_01v8__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_23=2.5575e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_23=-0.11838
.param sky130_fd_pr__pfet_01v8__ub_diff_23=2.6806e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_24=0.062257
.param sky130_fd_pr__pfet_01v8__ub_diff_24=2.5882e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_24=-0.016572
.param sky130_fd_pr__pfet_01v8__voff_diff_24=-0.007164
.param sky130_fd_pr__pfet_01v8__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_24=0.00061816
.param sky130_fd_pr__pfet_01v8__vsat_diff_24=-3126.4
.param sky130_fd_pr__pfet_01v8__vth0_diff_24=0.0093471
.param sky130_fd_pr__pfet_01v8__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_24=2.1916e-11
.param sky130_fd_pr__pfet_01v8__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_25=1.8662e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_25=0.14509
.param sky130_fd_pr__pfet_01v8__ub_diff_25=3.7411e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_25=-0.01248
.param sky130_fd_pr__pfet_01v8__voff_diff_25=-0.01901
.param sky130_fd_pr__pfet_01v8__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_25=0.00085089
.param sky130_fd_pr__pfet_01v8__vsat_diff_25=-21202.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_25=-0.020872
.param sky130_fd_pr__pfet_01v8__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_26=2.4441e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_26=0.35447
.param sky130_fd_pr__pfet_01v8__ub_diff_26=3.2678e-19
.param sky130_fd_pr__pfet_01v8__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_26=-0.018034
.param sky130_fd_pr__pfet_01v8__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_26=-0.0087068
.param sky130_fd_pr__pfet_01v8__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_26=0.0012768
.param sky130_fd_pr__pfet_01v8__vsat_diff_26=-7485.9
.param sky130_fd_pr__pfet_01v8__vth0_diff_26=-0.016578
.param sky130_fd_pr__pfet_01v8__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_27=-3.4302e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_27=-0.032055
.param sky130_fd_pr__pfet_01v8__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_27=0.017752
.param sky130_fd_pr__pfet_01v8__ub_diff_27=3.2461e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_27=-0.011438
.param sky130_fd_pr__pfet_01v8__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_27=-0.0078818
.param sky130_fd_pr__pfet_01v8__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_27=-0.027099
.param sky130_fd_pr__pfet_01v8__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_27=0.0011872
.param sky130_fd_pr__pfet_01v8__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_27=-0.010409
.param sky130_fd_pr__pfet_01v8__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_28=0.02972
.param sky130_fd_pr__pfet_01v8__ua_diff_28=-3.7577e-12
.param sky130_fd_pr__pfet_01v8__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_28=-0.011574
.param sky130_fd_pr__pfet_01v8__ub_diff_28=3.7012e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_28=-0.014576
.param sky130_fd_pr__pfet_01v8__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_28=-0.02451
.param sky130_fd_pr__pfet_01v8__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_28=0.014607
.param sky130_fd_pr__pfet_01v8__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_28=0.0015715
.param sky130_fd_pr__pfet_01v8__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_28=-0.0086025
.param sky130_fd_pr__pfet_01v8__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_29=0.058417
.param sky130_fd_pr__pfet_01v8__ua_diff_29=-6.6796e-13
.param sky130_fd_pr__pfet_01v8__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_29=-0.038418
.param sky130_fd_pr__pfet_01v8__ub_diff_29=4.1901e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_29=-0.013993
.param sky130_fd_pr__pfet_01v8__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_29=-0.026366
.param sky130_fd_pr__pfet_01v8__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_29=0.049839
.param sky130_fd_pr__pfet_01v8__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_29=0.0019461
.param sky130_fd_pr__pfet_01v8__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_29=-0.010094
.param sky130_fd_pr__pfet_01v8__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_30=-1.5243e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_30=0.07961
.param sky130_fd_pr__pfet_01v8__ub_diff_30=4.6877e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_30=-0.10304
.param sky130_fd_pr__pfet_01v8__k2_diff_30=-0.01506
.param sky130_fd_pr__pfet_01v8__voff_diff_30=-0.029429
.param sky130_fd_pr__pfet_01v8__a0_diff_30=0.12499
.param sky130_fd_pr__pfet_01v8__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_30=0.0021899
.param sky130_fd_pr__pfet_01v8__vth0_diff_30=-0.010409
.param sky130_fd_pr__pfet_01v8__u0_diff_31=0.00076283
.param sky130_fd_pr__pfet_01v8__vth0_diff_31=0.016967
.param sky130_fd_pr__pfet_01v8__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_31=1.8274e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_31=-0.075951
.param sky130_fd_pr__pfet_01v8__ub_diff_31=3.0138e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_31=-0.019051
.param sky130_fd_pr__pfet_01v8__voff_diff_31=-0.084009
.param sky130_fd_pr__pfet_01v8__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_31=-14746.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_32=-6821.2
.param sky130_fd_pr__pfet_01v8__u0_diff_32=0.00090881
.param sky130_fd_pr__pfet_01v8__vth0_diff_32=0.01388
.param sky130_fd_pr__pfet_01v8__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_32=2.73e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_32=-0.016583
.param sky130_fd_pr__pfet_01v8__ub_diff_32=3.457e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_32=-0.01911
.param sky130_fd_pr__pfet_01v8__voff_diff_32=0.009118
.param sky130_fd_pr__pfet_01v8__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_33=-0.001263
.param sky130_fd_pr__pfet_01v8__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_33=-20000.0
.param sky130_fd_pr__pfet_01v8__u0_diff_33=0.0010727
.param sky130_fd_pr__pfet_01v8__vth0_diff_33=-0.022734
.param sky130_fd_pr__pfet_01v8__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_33=6.2051e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_33=0.50111
.param sky130_fd_pr__pfet_01v8__ub_diff_33=3.5411e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_33=-0.016081
.param sky130_fd_pr__pfet_01v8__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_34=-0.01922
.param sky130_fd_pr__pfet_01v8__voff_diff_34=-0.060406
.param sky130_fd_pr__pfet_01v8__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_34=-11305.0
.param sky130_fd_pr__pfet_01v8__u0_diff_34=0.001349
.param sky130_fd_pr__pfet_01v8__vth0_diff_34=-0.0056167
.param sky130_fd_pr__pfet_01v8__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_34=5.1881e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_34=-0.37699
.param sky130_fd_pr__pfet_01v8__ub_diff_34=2.306e-19
.param sky130_fd_pr__pfet_01v8__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_35=-0.07957
.param sky130_fd_pr__pfet_01v8__ub_diff_35=-5.4359e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_35=0.0083879
.param sky130_fd_pr__pfet_01v8__voff_diff_35=0.00052667
.param sky130_fd_pr__pfet_01v8__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_35=-0.00048802
.param sky130_fd_pr__pfet_01v8__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_35=-0.031448
.param sky130_fd_pr__pfet_01v8__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_35=5.4688e-8
.param sky130_fd_pr__pfet_01v8__b1_diff_35=1.959e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_35=-5.4386e-12
.param sky130_fd_pr__pfet_01v8__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_36=-1.0533e-11
.param sky130_fd_pr__pfet_01v8__ua_diff_36=6.4807e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_36=1.1304
.param sky130_fd_pr__pfet_01v8__ub_diff_36=-5.9248e-21
.param sky130_fd_pr__pfet_01v8__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_36=0.014051
.param sky130_fd_pr__pfet_01v8__voff_diff_36=0.048748
.param sky130_fd_pr__pfet_01v8__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_36=-0.00029975
.param sky130_fd_pr__pfet_01v8__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_36=-0.0078078
.param sky130_fd_pr__pfet_01v8__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_36=-4.9985e-10
.param sky130_fd_pr__pfet_01v8__b0_diff_37=-2.4045e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_37=8.5392e-9
.param sky130_fd_pr__pfet_01v8__ua_diff_37=-6.2054e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_37=-0.044338
.param sky130_fd_pr__pfet_01v8__ub_diff_37=-2.5731e-21
.param sky130_fd_pr__pfet_01v8__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_37=0.0047513
.param sky130_fd_pr__pfet_01v8__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_37=-0.0091028
.param sky130_fd_pr__pfet_01v8__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_37=-0.00051198
.param sky130_fd_pr__pfet_01v8__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_37=-0.016784
.param sky130_fd_pr__pfet_01v8__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_38=-2.151e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_38=1.7904e-9
.param sky130_fd_pr__pfet_01v8__ua_diff_38=-2.9174e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_38=-0.013709
.param sky130_fd_pr__pfet_01v8__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_38=2.5002e-20
.param sky130_fd_pr__pfet_01v8__k2_diff_38=0.0034067
.param sky130_fd_pr__pfet_01v8__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_38=0.00018613
.param sky130_fd_pr__pfet_01v8__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_38=0.00026338
.param sky130_fd_pr__pfet_01v8__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_38=-0.019533
.param sky130_fd_pr__pfet_01v8__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_39=5.0e-10
.param sky130_fd_pr__pfet_01v8__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_39=8.2398e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_39=1.2806e-11
.param sky130_fd_pr__pfet_01v8__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_39=2.1839e-20
.param sky130_fd_pr__pfet_01v8__k2_diff_39=0.0071627
.param sky130_fd_pr__pfet_01v8__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_39=0.0063713
.param sky130_fd_pr__pfet_01v8__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_39=-8.9301e-5
.param sky130_fd_pr__pfet_01v8__vsat_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_39=-0.021886
.param sky130_fd_pr__pfet_01v8__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_40=-6.5314e-8
.param sky130_fd_pr__pfet_01v8__b1_diff_40=-1.198e-9
.param sky130_fd_pr__pfet_01v8__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_40=3.0902e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_40=-0.26607
.param sky130_fd_pr__pfet_01v8__ub_diff_40=2.7174e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_40=-0.031277
.param sky130_fd_pr__pfet_01v8__voff_diff_40=0.03868
.param sky130_fd_pr__pfet_01v8__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_40=20136.0
.param sky130_fd_pr__pfet_01v8__u0_diff_40=-0.00016379
.param sky130_fd_pr__pfet_01v8__vth0_diff_40=0.0026765
.param sky130_fd_pr__pfet_01v8__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_41=-7.0608e-8
.param sky130_fd_pr__pfet_01v8__b1_diff_41=3.4604e-10
.param sky130_fd_pr__pfet_01v8__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_41=-5.1088e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_41=0.032549
.param sky130_fd_pr__pfet_01v8__ub_diff_41=7.5534e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_41=-0.023281
.param sky130_fd_pr__pfet_01v8__voff_diff_41=-0.024626
.param sky130_fd_pr__pfet_01v8__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_41=20035.0
.param sky130_fd_pr__pfet_01v8__u0_diff_41=-4.5658e-5
.param sky130_fd_pr__pfet_01v8__vth0_diff_41=0.026137
.param sky130_fd_pr__pfet_01v8__u0_diff_42=0.00012907
.param sky130_fd_pr__pfet_01v8__vth0_diff_42=-0.047651
.param sky130_fd_pr__pfet_01v8__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_42=-6.299e-9
.param sky130_fd_pr__pfet_01v8__b1_diff_42=2.0752e-9
.param sky130_fd_pr__pfet_01v8__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_42=4.4904e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_42=0.042947
.param sky130_fd_pr__pfet_01v8__ub_diff_42=-1.7559e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_42=-0.0013346
.param sky130_fd_pr__pfet_01v8__voff_diff_42=-0.011769
.param sky130_fd_pr__pfet_01v8__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_42=20228.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_43=19828.0
.param sky130_fd_pr__pfet_01v8__u0_diff_43=-0.000155
.param sky130_fd_pr__pfet_01v8__vth0_diff_43=-0.034126
.param sky130_fd_pr__pfet_01v8__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_43=5.1711e-8
.param sky130_fd_pr__pfet_01v8__b1_diff_43=1.0663e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_43=-3.0557e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_43=-0.06169
.param sky130_fd_pr__pfet_01v8__ub_diff_43=1.0171e-21
.param sky130_fd_pr__pfet_01v8__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_43=0.0012972
.param sky130_fd_pr__pfet_01v8__voff_diff_43=-0.0049861
.param sky130_fd_pr__pfet_01v8__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_44=-0.040177
.param sky130_fd_pr__pfet_01v8__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_44=9.5149e-5
.param sky130_fd_pr__pfet_01v8__vth0_diff_44=-0.014011
.param sky130_fd_pr__pfet_01v8__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_44=-4.3729e-8
.param sky130_fd_pr__pfet_01v8__b1_diff_44=5.9219e-10
.param sky130_fd_pr__pfet_01v8__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_44=2.7637e-13
.param sky130_fd_pr__pfet_01v8__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_44=0.043802
.param sky130_fd_pr__pfet_01v8__ub_diff_44=7.4297e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_44=-0.0060597
.param sky130_fd_pr__pfet_01v8__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_45=0.0036376
.param sky130_fd_pr__pfet_01v8__voff_diff_45=-0.0089003
.param sky130_fd_pr__pfet_01v8__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_45=20022.0
.param sky130_fd_pr__pfet_01v8__u0_diff_45=-3.1766e-5
.param sky130_fd_pr__pfet_01v8__vth0_diff_45=-0.0090051
.param sky130_fd_pr__pfet_01v8__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_45=-1.2637e-8
.param sky130_fd_pr__pfet_01v8__b1_diff_45=5.0054e-10
.param sky130_fd_pr__pfet_01v8__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_45=-9.1068e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_45=0.003075
.param sky130_fd_pr__pfet_01v8__ub_diff_45=8.5731e-21
.param sky130_fd_pr__pfet_01v8__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_46=-0.020789
.param sky130_fd_pr__pfet_01v8__ub_diff_46=-1.0587e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_46=0.0037416
.param sky130_fd_pr__pfet_01v8__voff_diff_46=-0.0015691
.param sky130_fd_pr__pfet_01v8__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_46=-0.00043944
.param sky130_fd_pr__pfet_01v8__vsat_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_46=-0.0074705
.param sky130_fd_pr__pfet_01v8__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_46=3.1294e-9
.param sky130_fd_pr__pfet_01v8__b1_diff_46=2.2449e-9
.param sky130_fd_pr__pfet_01v8__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_46=1.9375e-12
.param sky130_fd_pr__pfet_01v8__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_47=4.76e-10
.param sky130_fd_pr__pfet_01v8__ua_diff_47=5.6931e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_47=-0.022087
.param sky130_fd_pr__pfet_01v8__ub_diff_47=1.5369e-20
.param sky130_fd_pr__pfet_01v8__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_47=-0.026507
.param sky130_fd_pr__pfet_01v8__voff_diff_47=0.0055712
.param sky130_fd_pr__pfet_01v8__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_47=-0.00040161
.param sky130_fd_pr__pfet_01v8__vsat_diff_47=19939.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_47=0.04187
.param sky130_fd_pr__pfet_01v8__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_47=-1.1127e-7
.param sky130_fd_pr__pfet_01v8__b0_diff_48=-7.0103e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_48=-1.7236e-10
.param sky130_fd_pr__pfet_01v8__ua_diff_48=8.7575e-12
.param sky130_fd_pr__pfet_01v8__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_48=0.0069841
.param sky130_fd_pr__pfet_01v8__ub_diff_48=1.0058e-19
.param sky130_fd_pr__pfet_01v8__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_48=-0.017287
.param sky130_fd_pr__pfet_01v8__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_48=-0.028186
.param sky130_fd_pr__pfet_01v8__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_48=0.00044832
.param sky130_fd_pr__pfet_01v8__vsat_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_48=-0.024556
.param sky130_fd_pr__pfet_01v8__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_49=5.7731e-8
.param sky130_fd_pr__pfet_01v8__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_49=1.4765e-8
.param sky130_fd_pr__pfet_01v8__ua_diff_49=6.0464e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_49=-0.98866
.param sky130_fd_pr__pfet_01v8__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__ub_diff_49=-1.3903e-19
.param sky130_fd_pr__pfet_01v8__k2_diff_49=-0.011802
.param sky130_fd_pr__pfet_01v8__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__voff_diff_49=0.0021743
.param sky130_fd_pr__pfet_01v8__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__u0_diff_49=-0.00012869
.param sky130_fd_pr__pfet_01v8__vsat_diff_49=20208.0
.param sky130_fd_pr__pfet_01v8__vth0_diff_49=-0.026247
.param sky130_fd_pr__pfet_01v8__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_50=3.6372e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_50=-0.77531
.param sky130_fd_pr__pfet_01v8__ub_diff_50=1.5241e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_50=-0.037862
.param sky130_fd_pr__pfet_01v8__voff_diff_50=0.027312
.param sky130_fd_pr__pfet_01v8__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_50=90.881
.param sky130_fd_pr__pfet_01v8__u0_diff_50=0.00046495
.param sky130_fd_pr__pfet_01v8__vth0_diff_50=-0.023191
.param sky130_fd_pr__pfet_01v8__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__kt1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__agidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__ua_diff_51=2.1342e-11
.param sky130_fd_pr__pfet_01v8__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__nfactor_diff_51=-0.19662
.param sky130_fd_pr__pfet_01v8__ub_diff_51=2.8241e-19
.param sky130_fd_pr__pfet_01v8__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__ags_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__k2_diff_51=-0.036739
.param sky130_fd_pr__pfet_01v8__voff_diff_51=0.052482
.param sky130_fd_pr__pfet_01v8__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__vsat_diff_51=89.681
.param sky130_fd_pr__pfet_01v8__u0_diff_51=0.00082673
.param sky130_fd_pr__pfet_01v8__vth0_diff_51=0.02896
.param sky130_fd_pr__pfet_01v8__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8__keta_diff_51=0.0
.include "sky130_fd_pr__pfet_01v8.pm3.spice"