* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre=0.0
.subckt sky130_fd_pr__pfet_01v8_hvt d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__pfet_01v8_hvt d g s b sky130_fd_pr__pfet_01v8_hvt__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos lmin=2.0e-05 lmax=0.0001 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.1096107+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43657182 k2=0.027786788 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.62938688+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='7.7456776+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.019607098 ua=-2.7648397e-10 ub=2.34385173e-18 uc=-7.7670696e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=200000.0 a0=1.5015529 ags=0.3818821 a1=0.0 a2=1.0 b0=0.0 b1=0.0 keta=-0.013169082 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.075489662 pdiblc1=0.39 pdiblc2=0.0036275994 pdiblcb=-9.5744039e-5 drout=0.56 pscbe1=746475130.0 pscbe2=9.5049925e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.7923891 agidl=6.8812e-10 bgidl=1154444600.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.44169 kt2=-0.037961 at=0.0 ute=-0.30066 ua1=2.2116e-9 ub1=-7.9359e-19 uc1=1.1985e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.1096107+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43657182 k2=0.027786788 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.62938688+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='7.7456776+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.019607098 ua=-2.7648397e-10 ub=2.34385173e-18 uc=-7.7670696e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=200000.0 a0=1.5015529 ags=0.3818821 a1=0.0 a2=1.0 b0=0.0 b1=0.0 keta=-0.013169082 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.075489662 pdiblc1=0.39 pdiblc2=0.0036275994 pdiblcb=-9.5744039e-5 drout=0.56 pscbe1=746475130.0 pscbe2=9.5049925e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.7923891 agidl=6.8812e-10 bgidl=1154444600.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.44169 kt2=-0.037961 at=0.0 ute=-0.30066 ua1=2.2116e-9 ub1=-7.9359e-19 uc1=1.1985e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108727938e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.052274411e-09 wvth0=-8.831651785e-08 pvth0=7.055491799e-13 k1=4.360518078e-01 lk1=4.154309705e-09 wk1=5.202494200e-08 pk1=-4.156204984e-13 k2=2.819103967e-02 lk2=-3.229514006e-09 wk2=-4.044360936e-08 pk2=3.230987375e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.285207292e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-6.919566331e-09 wvoff=-8.665459790e-08 pvoff=6.922723176e-13 nfactor='7.724686277e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.676969498e-07 wnfactor=2.100089957e-06 pnfactor=-1.677734565e-11 eta0=0.08 etab=-0.07 u0=1.932456476e-02 lu0=2.257121325e-09 wu0=2.826621373e-08 pu0=-2.258151068e-13 ua=-3.021630050e-10 lua=2.051464722e-16 wua=2.569075027e-15 pua=-2.052400641e-20 ub=2.324401486e-18 lub=1.553854689e-25 wub=1.945911736e-24 pub=-1.554563589e-29 uc=-7.712273168e-11 luc=-4.377615734e-18 wuc=-5.482143144e-17 puc=4.379612890e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.943880576e+05 lvsat=4.483307809e-02 wvsat=5.614502657e-01 pvsat=-4.485353184e-6 a0=1.524414571e+00 la0=-1.826389211e-07 wa0=-2.287210140e-06 pa0=1.827222447e-11 ags=4.009303173e-01 lags=-1.521737318e-07 wags=-1.905690749e-06 pags=1.522431565e-11 a1=0.0 a2=9.848810403e-01 la2=1.207035148e-07 wa2=1.511585270e-06 pa2=-1.207585822e-11 b0=0.0 b1=0.0 keta=-1.635811733e-02 lketa=2.547678869e-08 wketa=3.190490233e-07 pketa=-2.548841171e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.175946087e-01 lpclm=-3.363709457e-07 wpclm=-4.212415583e-06 ppclm=3.365244048e-11 pdiblc1=0.39 pdiblc2=3.389656634e-03 lpdiblc2=1.900893826e-09 wpdiblc2=2.380513203e-08 ppdiblc2=-1.901761051e-13 pdiblcb=-1.467644794e-04 lpdiblcb=4.075956659e-10 wpdiblcb=5.104371697e-09 ppdiblcb=-4.077816192e-14 drout=0.56 pscbe1=7.505188577e+08 lpscbe1=-3.230481493e+01 wpscbe1=-4.045572532e+02 ppscbe1=3.231955303e-3 pscbe2=9.463108264e-09 lpscbe2=3.346077183e-16 wpscbe2=4.190334466e-15 ppscbe2=-3.347603731e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.831979289e+00 lbeta0=-3.162808702e-07 wbeta0=-3.960825046e-06 pbeta0=3.164251638e-11 agidl=6.551754237e-10 lagidl=2.631899371e-16 wagidl=3.295960625e-15 pagidl=-2.633100096e-20 bgidl=1.142776530e+09 lbgidl=9.321469104e+01 wbgidl=1.167339279e+03 pbgidl=-9.325721745e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.425036582e-01 lkt1=6.500209282e-09 wkt1=8.140293693e-08 pkt1=-6.503174808e-13 kt2=-3.814118335e-02 lkt2=1.439461387e-09 wkt2=1.802655567e-08 pkt2=-1.440118098e-13 at=1.983225665e+04 lat=-1.584373202e-01 wat=-1.984130453e+00 pat=1.585096025e-5 ute=-3.004779279e-01 lute=-1.454550081e-09 wute=-1.821551328e-08 pute=1.455213676e-13 ua1=2.227223445e-09 lua1=-1.248136750e-16 wua1=-1.563057322e-15 pua1=1.248706175e-20 ub1=-8.067528284e-19 lub1=1.051561247e-25 wub1=1.316883352e-24 pub1=-1.052040991e-29 uc1=1.211396142e-10 luc1=-1.030256012e-17 wuc1=-1.290202538e-16 puc1=1.030726035e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.122594846e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.826102235e-08 wvth0=1.365094275e-07 pvth0=-1.912522886e-13 k1=4.493657172e-01 lk1=-4.895314383e-08 wk1=-5.951765964e-07 pk1=2.165982302e-12 k2=1.965123111e-02 lk2=3.083467214e-08 wk2=2.815734565e-07 pk2=-9.613854759e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=5.442199869e-01 ldsub=6.294442095e-08 wdsub=1.578721228e-06 pdsub=-6.297313746e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.377410065e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.985892130e-08 wvoff=-3.048281824e-07 pvoff=1.562538384e-12 nfactor='8.043758479e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.105040586e-06 wnfactor=-2.178506005e-06 pnfactor=2.894174196e-13 eta0=7.401064685e-02 leta0=2.389075108e-08 weta0=5.992085608e-07 peta0=-2.390165052e-12 etab=-6.476402461e-02 letab=-2.088562516e-08 wetab=-5.238364148e-07 petab=2.089515360e-12 u0=2.365925872e-02 lu0=-1.503340935e-08 wu0=-3.333684774e-08 pu0=1.991149696e-14 ua=9.272450516e-11 lua=-1.370008470e-15 wua=-3.121327775e-15 pua=2.174270613e-21 ub=2.623200850e-18 lub=-1.036486351e-24 wub=-2.333901187e-24 pub=1.525981486e-30 uc=-8.615807197e-11 luc=3.166318211e-17 wuc=1.275182190e-16 puc=-2.893678725e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.799149686e+05 lvsat=-2.963226514e-01 wvsat=-6.048539334e-01 pvsat=1.668826468e-7 a0=1.152376958e+00 la0=1.301370755e-06 wa0=4.827307396e-06 pa0=-1.010666109e-11 ags=1.060806321e-01 lags=1.023943332e-06 wags=2.508397131e-06 pags=-2.382907068e-12 a1=0.0 a2=1.229084975e+00 la2=-8.533942343e-07 wa2=-3.023170540e-06 pa2=6.012693192e-12 b0=0.0 b1=0.0 keta=3.501192289e-02 lketa=-1.794316236e-07 wketa=-6.207023588e-07 pketa=1.199704925e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.647293317e-01 lpclm=2.385330551e-06 wpclm=8.603689119e-06 ppclm=-1.746933508e-11 pdiblc1=0.39 pdiblc2=7.217847004e-03 lpdiblc2=-1.336925990e-08 wpdiblc2=-4.584503763e-08 ppdiblc2=8.764936711e-14 pdiblcb=6.199588191e-04 lpdiblcb=-2.650763898e-09 wpdiblcb=-4.414829700e-09 ppdiblcb=-2.807305045e-15 drout=0.56 pscbe1=6.851606705e+08 lpscbe1=2.284004973e+02 wpscbe1=8.091145064e+02 ppscbe1=-1.609223568e-3 pscbe2=1.011912642e-08 lpscbe2=-2.282163411e-15 wpscbe2=-6.284641909e-15 ppscbe2=8.307281707e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.340918808e+00 lbeta0=1.642495549e-06 wbeta0=-6.968142227e-06 pbeta0=4.363831367e-11 agidl=1.187654568e-09 lagidl=-1.860800146e-15 wagidl=-6.591992552e-15 pagidl=1.311075883e-20 bgidl=1.331365855e+09 lbgidl=-6.590436080e+02 wbgidl=-2.334678558e+03 pbgidl=4.643372143e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.277110086e-01 lkt1=-5.250574678e-08 wkt1=-3.270417800e-07 pkt1=9.789153974e-13 kt2=-3.548113669e-02 lkt2=-9.171118947e-09 wkt2=-1.081851686e-08 pkt2=-2.895256535e-14 at=-3.136423608e+05 lat=1.171749577e+00 wat=5.261722303e+00 pat=-1.305180443e-5 ute=-2.935034937e-01 lute=-2.927466138e-08 wute=-9.557452919e-07 pute=3.885205776e-12 ua1=1.930766960e-09 lua1=1.057712705e-15 wua1=7.521818200e-15 pua1=-2.375132567e-20 ub1=-5.690430214e-19 lub1=-8.430373928e-25 wub1=-5.130996646e-24 pub1=1.519934518e-29 uc1=8.453246673e-11 luc1=1.357185922e-16 wuc1=1.835089605e-15 puc1=-6.803852856e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.096737981e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.164922517e-09 wvth0=-1.188561471e-07 pvth0=3.166366418e-13 k1=4.209874975e-01 lk1=7.487445918e-09 wk1=8.705142160e-07 pk1=-7.490861840e-13 k2=3.664638724e-02 lk2=-2.966484037e-09 wk2=-3.510315989e-07 pk2=2.967837406e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=6.245231430e-01 ldsub=-9.676811721e-08 wdsub=-6.455257977e-06 pdsub=9.681226476e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.223681671e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.156578288e-10 wvoff=4.448135493e-07 pvoff=7.159843262e-14 nfactor='7.352043218e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.706911459e-07 wnfactor=1.158352041e-05 pnfactor=-2.708146407e-11 eta0=1.024505933e-01 leta0=-3.267260519e-08 weta0=-2.246083570e-06 peta0=3.268751109e-12 etab=-7.530273474e-02 letab=7.449926597e-11 wetab=5.305153957e-07 petab=-7.453325403e-15 u0=1.600429451e-02 lu0=1.913193151e-10 wu0=-1.370149861e-08 pu0=-1.914065988e-14 ua=-5.894234371e-10 lua=-1.330489245e-17 wua=-2.697381327e-15 pua=1.331096241e-21 ub=2.074848117e-18 lub=5.411594944e-26 wub=1.155540208e-24 pub=-5.414063822e-30 uc=-6.957681104e-11 luc=-1.314790313e-18 wuc=-8.411295202e-17 puc=1.315390146e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.333042000e+05 lvsat=-4.732892029e-03 wvsat=-7.590231250e-01 pvsat=4.735051269e-7 a0=1.807850106e+00 la0=-2.280124534e-09 wa0=-3.689988340e-07 pa0=2.281164773e-13 ags=6.297427835e-01 lags=-1.755261114e-08 wags=4.273315173e-07 pags=1.756061899e-12 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-5.402520275e-02 lketa=-2.348355581e-09 wketa=-1.356217703e-07 pketa=2.349426948e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.430702329e-01 lpclm=-1.682576948e-08 wpclm=-1.026241271e-06 ppclm=1.683344573e-12 pdiblc1=3.865953011e-01 lpdiblc1=6.771503502e-09 wpdiblc1=3.406252192e-07 ppdiblc1=-6.774592797e-13 pdiblc2=5.097534716e-04 lpdiblc2=-2.773391177e-11 wpdiblc2=-3.170196810e-09 ppdiblc2=2.774656454e-15 pdiblcb=-6.978912554e-04 lpdiblcb=-2.973142036e-11 wpdiblcb=-7.321909342e-09 ppdiblcb=2.974498443e-15 drout=5.816813724e-01 ldrout=-4.312143120e-08 wdrout=-2.169126392e-06 pdrout=4.314110406e-12 pscbe1=800000000.0 pscbe2=9.004001941e-09 lpscbe2=-6.432579521e-17 wpscbe2=-5.343520813e-15 ppscbe2=6.435514193e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.280633849e+00 lbeta0=-2.264755038e-07 wbeta0=3.580778026e-06 pbeta0=2.265788264e-11 agidl=2.761605116e-10 lagidl=-4.795696251e-17 wagidl=-2.412295192e-15 pagidl=4.797884144e-21 bgidl=1.009479675e+09 lbgidl=-1.885384214e+01 wbgidl=-9.484000280e+02 pbgidl=1.886244364e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.571230211e-01 lkt1=5.990922543e-09 wkt1=4.665148474e-07 pkt1=-5.993655721e-13 kt2=-4.035397695e-02 lkt2=5.203268623e-10 wkt2=7.980590052e-10 pkt2=-5.205642458e-14 at=2.796698942e+05 lat=-8.271367424e-03 wat=-1.716772285e+00 pat=8.275140987e-7 ute=-4.014196268e-01 lute=1.853564981e-07 wute=1.032166948e-05 pute=-1.854410615e-11 ua1=2.276780712e-09 lua1=3.695363340e-16 wua1=1.416838973e-14 pua1=-3.697049238e-20 ub1=-8.879763809e-19 lub1=-2.087204022e-25 wub1=-7.988004532e-24 pub1=2.088156246e-29 uc1=1.581711189e-10 luc1=-1.073911389e-17 wuc1=-2.126081405e-15 puc1=1.074401329e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.104347290e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.359695254e-09 wvth0=1.216943736e-07 pvth0=7.876344834e-14 k1=3.626009089e-01 lk1=6.522419181e-08 wk1=3.379529178e-07 pk1=-2.224522931e-13 k2=6.088486525e-02 lk2=-2.693518778e-08 wk2=-1.714622965e-07 pk2=1.192130445e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=7.469753064e-01 ldsub=-2.178573881e-07 wdsub=1.782716347e-06 pdsub=1.534940806e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.869161829e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.311393861e-08 wvoff=6.972527454e-07 pvoff=-1.780311152e-13 nfactor='7.850860776e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.225745730e-07 wnfactor=-1.208353807e-05 pnfactor=-3.677819941e-12 eta0=1.378002277e-01 leta0=-6.762879820e-08 weta0=1.993919478e-06 peta0=-9.240607050e-13 etab=-1.483283986e-01 letab=7.228738745e-08 wetab=1.038020206e-06 petab=-5.093096073e-13 u0=1.923746476e-02 lu0=-3.005865755e-09 wu0=-3.613183911e-08 pu0=3.040030940e-15 ua=-3.329492658e-10 lua=-2.669245063e-16 wua=-2.182009776e-15 pua=8.214607756e-22 ub=2.323395052e-18 lub=-1.916646575e-25 wub=-3.491645699e-24 pub=-8.186010938e-31 uc=-6.477667493e-11 luc=-6.061500909e-18 wuc=-3.323576763e-16 puc=3.770207751e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.983985711e+05 lvsat=-6.910276280e-02 wvsat=-5.481775556e-01 pvsat=2.650062686e-7 a0=1.788834346e+00 la0=1.652398926e-08 wa0=4.815434942e-06 pa0=-4.898614551e-12 ags=4.309367551e-01 lags=1.790407062e-07 wags=3.406763338e-06 pags=-1.190208846e-12 a1=0.0 a2=8.148138538e-01 la2=-1.464897560e-08 wa2=-1.482061217e-06 pa2=1.465565876e-12 b0=0.0 b1=0.0 keta=-5.314527244e-02 lketa=-3.218492269e-09 wketa=2.107756890e-09 pketa=9.874609720e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.633949386e-01 lpclm=-3.692426118e-08 wpclm=-7.384055170e-07 ppclm=1.398712431e-12 pdiblc1=3.720535046e-01 lpdiblc1=2.115144982e-08 wpdiblc1=1.795468297e-06 ppdiblc1=-2.116109954e-12 pdiblc2=7.537206750e-04 lpdiblc2=-2.689857602e-10 wpdiblc2=-4.668789910e-09 ppdiblc2=4.256570213e-15 pdiblcb=-1.671969296e-03 lpdiblcb=9.335051313e-10 wpdiblcb=1.653242344e-07 ppdiblcb=-1.677500937e-13 drout=5.457651998e-01 ldrout=-7.605005539e-09 wdrout=1.424129443e-06 pdrout=7.608475095e-13 pscbe1=7.969604563e+08 lpscbe1=3.005713570e+00 wpscbe1=3.040930392e+02 ppscbe1=-3.007084837e-4 pscbe2=9.233762175e-09 lpscbe2=-2.915287980e-16 wpscbe2=-1.127610960e-15 ppscbe2=2.266527416e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=2.992863204e+00 lbeta0=2.035832253e-06 wbeta0=3.922123529e-05 pbeta0=-1.258589633e-11 agidl=2.412136287e-10 lagidl=-1.339903841e-17 wagidl=1.083062081e-15 pagidl=1.341430196e-21 bgidl=9.935672924e+08 lbgidl=-3.118563934e+00 wbgidl=6.435642293e+02 pbgidl=3.119986685e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.754280130e-01 lkt1=2.409217992e-08 wkt1=1.663817167e-07 pkt1=-3.025729233e-13 kt2=-3.523070398e-02 lkt2=-4.545924082e-09 wkt2=-1.842662778e-07 pkt2=1.309481461e-13 at=4.439247213e+05 lat=-1.706980384e-01 wat=-1.363097581e+00 pat=4.777757946e-7 ute=-2.560929686e-01 lute=4.164732565e-08 wute=-1.709417433e-05 pute=8.566599321e-12 ua1=3.501774071e-09 lua1=-8.418228484e-16 wua1=-5.133902149e-14 pua1=2.780782134e-20 ub1=-1.658531144e-18 lub1=5.532580868e-25 wub1=3.669336537e-23 pub1=-2.330250380e-29 uc1=3.529363748e-10 luc1=-2.033366325e-16 wuc1=-1.144416457e-15 puc1=1.036623125e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.095738847e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.512856226e-10 wvth0=3.137677521e-07 pvth0=-1.513546421e-14 k1=5.154033531e-01 lk1=-9.476339101e-09 wk1=-2.056382044e-06 pk1=9.480662397e-13 k2=-7.801580673e-04 lk2=3.210992167e-09 wk2=7.295108724e-07 pk2=-3.212457086e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.784316906e-01 ldsub=1.119952944e-08 wdsub=7.214435814e-06 pdsub=-1.120463889e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.487571068e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.427888935e-09 wvoff=-5.730686445e-07 pvoff=4.429909027e-13 nfactor='7.298367773e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.752268156e-08 wnfactor=-9.881283289e-06 pnfactor=-4.754436236e-12 eta0=3.390588200e-02 leta0=-1.683796940e-08 weta0=-3.342112243e-06 peta0=1.684565122e-12 etab=-4.349753485e-04 letab=-1.327035823e-11 wetab=-6.505431706e-09 petab=1.327641243e-15 u0=1.283424712e-02 lu0=1.244752524e-10 wu0=-4.439906714e-09 pu0=-1.245320405e-14 ua=-9.427720475e-10 lua=3.119955704e-17 wua=5.883201561e-15 pua=-3.121379091e-21 ub=1.974182722e-18 lub=-2.094522568e-26 wub=-9.452492600e-24 pub=2.095478131e-30 uc=-7.609646532e-11 luc=-5.275949820e-19 wuc=3.308804176e-16 puc=5.278356814e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.803911417e+04 lvsat=-4.852350721e-04 wvsat=-1.054000810e-01 pvsat=4.854564460e-8 a0=1.800777597e+00 la0=1.068529245e-08 wa0=-3.018135991e-06 pa0=-1.069016729e-12 ags=8.964161366e-01 lags=-4.851819906e-08 wags=-8.956937133e-06 pags=4.854033404e-12 a1=0.0 a2=7.703722924e-01 la2=7.077170512e-09 wa2=2.964122434e-06 pa2=-7.080399259e-13 b0=0.0 b1=0.0 keta=-6.383587559e-02 lketa=2.007822894e-09 wketa=6.149905017e-07 pketa=-2.008738903e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.757783535e-01 lpclm=5.908858790e-09 wpclm=3.331936055e-06 ppclm=-5.911554530e-13 pdiblc1=4.384124393e-01 lpdiblc1=-1.128944260e-08 wpdiblc1=-4.843452603e-06 ppdiblc1=1.129459307e-12 pdiblc2=7.604466525e-04 lpdiblc2=-2.722738888e-10 wpdiblc2=-5.168177975e-08 ppdiblc2=2.723981056e-14 pdiblcb=2.375467952e-04 wpdiblcb=-1.778142149e-7 drout=5.018998453e-01 ldrout=1.383945029e-08 wdrout=5.812666112e-06 pdrout=-1.384576412e-12 pscbe1=8.060790874e+08 lpscbe1=-1.452111603e+00 wpscbe1=-6.081860784e+02 ppscbe1=1.452774086e-4 pscbe2=8.048535097e-09 lpscbe2=2.878931638e-16 wpscbe2=6.242502687e-14 ppscbe2=-2.880245064e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.235084956e-09 lalpha0=-5.549089824e-16 walpha0=-1.135602804e-13 palpha0=5.551621430e-20 alpha1=9.276134311e-11 lalpha1=3.538762194e-18 walpha1=7.241959311e-16 palpha1=-3.540376648e-22 beta0=7.705846421e+00 lbeta0=-2.682038519e-07 wbeta0=-4.141066586e-05 pbeta0=2.683262118e-11 agidl=2.471771017e-10 lagidl=-1.631440147e-17 wagidl=4.883145081e-16 pagidl=1.632184442e-21 bgidl=9.924854795e+08 lbgidl=-2.589698023e+00 wbgidl=7.517948818e+02 pbgidl=2.590879495e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.266178953e-01 lkt1=2.303776654e-10 wkt1=-4.053953333e-07 pkt1=-2.304827683e-14 kt2=-4.494262190e-02 lkt2=2.019412340e-10 wkt2=1.249191549e-07 pkt2=-2.020333636e-14 at=9.513885628e+04 lat=-1.870925171e-04 wat=-4.240790133e-01 pat=1.871778724e-8 ute=-1.665587714e-01 lute=-2.123257317e-09 wute=-5.425330174e-09 pute=2.124225989e-13 ua1=1.681101245e-09 lua1=4.824947608e-17 wua1=1.541690583e-14 pua1=-4.827148846e-21 ub1=-4.297318726e-19 lub1=-4.746501319e-26 wub1=-2.068624591e-23 pub1=4.748666767e-30 uc1=-5.422306194e-11 luc1=-4.288598690e-18 wuc1=-1.810019196e-15 puc1=4.290555235e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.111883068e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.007655793e-09 wvth0=1.928926426e-06 pvth0=-4.009484166e-13 k1=5.190311829e-01 lk1=-1.034291882e-08 wk1=-2.419330537e-06 pk1=1.034763746e-12 k2=-2.503657329e-03 lk2=3.622684435e-09 wk2=9.019394281e-07 pk2=-3.624337176e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.036552333e-01 ldsub=5.174381798e-09 wdsub=4.690930795e-06 pdsub=-5.176742454e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.671694757e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.972639033e-11 wvoff=1.269008249e-06 pvoff=2.973995211e-15 nfactor='7.513625325e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.895889874e-09 wnfactor=-3.141685896e-05 pnfactor=3.897667257e-13 eta0=-3.658421472e-02 weta0=3.710113328e-6 etab=-4.905300834e-04 letab=1.309705708e-18 wetab=-9.474236925e-10 petab=-1.310303216e-22 u0=1.302198035e-02 lu0=7.963141643e-11 wu0=-2.322179421e-08 pu0=-7.966774587e-15 ua=-8.720118943e-10 lua=1.429707924e-17 wua=-1.196041982e-15 pua=-1.430360186e-21 ub=1.900026297e-18 lub=-3.231480537e-27 wub=-2.033466978e-24 pub=3.232954803e-31 uc=-8.030829580e-11 luc=4.784849643e-19 wuc=7.522556176e-16 puc=-4.787032587e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.633349567e+04 lvsat=-7.781398148e-05 wvsat=6.523958257e-02 pvsat=7.784948178e-9 a0=1.813161022e+00 la0=7.727263646e-09 wa0=-4.257043477e-06 pa0=-7.730788978e-13 ags=5.002652128e-01 lags=4.611037211e-08 wags=3.067622845e-05 pags=-4.613140858e-12 a1=0.0 a2=7.862174314e-01 la2=3.292242150e-09 wa2=1.378885644e-06 pa2=-3.293744137e-13 b0=0.0 b1=0.0 keta=-5.556141279e-02 lketa=3.130196629e-11 wketa=-2.128332752e-07 pketa=-3.131624688e-15 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.970489189e-01 lpclm=8.279588369e-10 wpclm=1.203909110e-06 ppclm=-8.283365683e-14 pdiblc1=3.971394206e-01 lpdiblc1=-1.430556614e-09 wpdiblc1=-7.142677733e-07 ppdiblc1=1.431209262e-13 pdiblc2=-2.576915399e-04 lpdiblc2=-2.907121879e-11 wpdiblc2=5.017848898e-08 ppdiblc2=2.908448166e-15 pdiblcb=-2.724839315e-02 lpdiblcb=6.565566475e-09 wpdiblcb=2.572033743e-06 ppdiblcb=-6.568561818e-13 drout=5.640284291e-01 ldrout=-1.001204524e-09 wdrout=-4.030266976e-07 pdrout=1.001661294e-13 pscbe1=7.999813105e+08 lpscbe1=4.464350172e-03 wpscbe1=1.869798174e+00 ppscbe1=-4.466386898e-7 pscbe2=1.076745325e-08 lpscbe2=-3.615748147e-16 wpscbe2=-2.095908306e-13 ppscbe2=3.617397723e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-1.319903354e-09 lalpha0=5.540107511e-17 walpha0=1.420551142e-13 palpha0=-5.542635018e-21 alpha1=1.075759376e-10 walpha1=-7.579393929e-16 beta0=6.498208410e+00 lbeta0=2.026463977e-08 wbeta0=7.940823008e-05 pbeta0=-2.027388490e-12 agidl=-2.545138795e-11 lagidl=4.880836585e-17 wagidl=2.776360133e-14 pagidl=-4.883063321e-21 bgidl=1.009965861e+09 lbgidl=-6.765236785e+00 wbgidl=-9.970407720e+02 pbgidl=6.768323221e-4 cgidl=2.541335236e+02 lcgidl=1.095612521e-05 wcgidl=4.588740156e-03 pcgidl=-1.096112361e-9 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.015072196e-01 lkt1=-5.767809451e-09 wkt1=-2.917608508e-06 pkt1=5.770440842e-13 kt2=-4.678647856e-02 lkt2=6.423832743e-10 wkt2=3.093889413e-07 pkt2=-6.426763424e-14 at=9.211512097e+04 lat=5.351871368e-04 wat=-1.215675333e-01 pat=-5.354312999e-8 ute=-1.968199601e-01 lute=5.105232829e-09 wute=3.022074116e-06 pute=-5.107561938e-13 ua1=1.732232133e-09 lua1=3.603584080e-17 wua1=1.030148431e-14 pua1=-3.605228107e-21 ub1=-4.797891031e-19 lub1=-3.550784255e-26 wub1=-1.567823916e-23 pub1=3.552404194e-30 uc1=-6.033673320e-11 luc1=-2.828226037e-18 wuc1=-1.198373152e-15 puc1=2.829516330e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.095735939e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.409836289e-09 wvth0=3.134768862e-07 pvth0=-1.410479485e-13 k1=4.964210488e-01 lk1=-7.181586072e-09 wk1=-1.572856055e-07 pk1=7.184862455e-13 k2=-7.401941116e-03 lk2=4.897821019e-09 wk2=1.391991276e-06 pk2=-4.900055503e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.336286821e-01 ldsub=1.871111750e-08 wdsub=1.169678066e-05 pdsub=-1.871965389e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.487048067e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.464746941e-09 wvoff=-5.783010426e-07 pvoff=3.466327627e-13 nfactor='7.034567078e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=8.475447048e-08 wnfactor=1.651082129e-05 pnfactor=-8.479313716e-12 eta0=-1.428617406e-01 leta0=1.975380374e-08 weta0=1.434271451e-05 peta0=-1.976281582e-12 etab=-1.435743743e-02 letab=2.577442070e-09 wetab=1.386375947e-06 petab=-2.578617951e-13 u0=1.375183258e-02 lu0=-4.800979094e-11 wu0=-9.624031490e-08 pu0=4.803169397e-15 ua=-6.974822802e-10 lua=-1.670346527e-17 wua=-1.865696578e-14 pua=1.671108572e-21 ub=1.792656427e-18 lub=1.640004684e-26 wub=8.708418478e-24 pub=-1.640752887e-30 uc=-7.907655520e-11 luc=2.977100152e-19 wuc=6.290253630e-16 puc=-2.978458364e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.984818477e+04 lvsat=1.119777288e-03 wvsat=7.140665456e-01 pvsat=-1.120288153e-7 a0=1.854219846e+00 la0=8.735570988e-10 wa0=-8.364799074e-06 pa0=-8.739556330e-14 ags=7.733176917e-01 wags=3.358523358e-6 a1=0.0 a2=8.290347267e-01 la2=-4.334781278e-09 wa2=-2.904797287e-06 pa2=4.336758892e-13 b0=8.294764088e-25 lb0=-1.541747801e-31 wb0=-8.298548325e-29 pb0=1.542451177e-35 b1=0.0 keta=-2.919241805e-02 lketa=-4.866751944e-09 wketa=-2.850935756e-06 pketa=4.868972254e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.722944029e-01 lpclm=5.512430626e-09 wpclm=3.680490053e-06 ppclm=-5.514945507e-13 pdiblc1=2.985345433e-01 lpdiblc1=1.675311901e-08 wpdiblc1=9.150718511e-06 ppdiblc1=-1.676076212e-12 pdiblc2=-2.508230397e-03 lpdiblc2=3.863098635e-10 wpdiblc2=2.753350487e-07 ppdiblc2=-3.864861058e-14 pdiblcb=1.424476603e-02 lpdiblcb=-4.858170014e-10 wpdiblcb=-1.579175176e-06 ppdiblcb=4.860386408e-14 drout=7.214186447e-01 ldrout=-3.035611431e-08 wdrout=-1.614922871e-05 pdrout=3.036996337e-12 pscbe1=8.000479988e+08 lpscbe1=-7.481570262e-03 wpscbe1=-4.802068072e+00 ppscbe1=7.484983504e-7 pscbe2=8.717893628e-09 lpscbe2=-1.702259894e-17 wpscbe2=-4.541363702e-15 ppscbe2=1.703036499e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-4.486325314e-09 lalpha0=6.495211042e-16 walpha0=4.588417687e-13 palpha0=-6.498174287e-20 alpha1=1.075759376e-10 walpha1=-7.579393929e-16 beta0=5.698187331e+00 lbeta0=1.710045819e-07 wbeta0=1.594468366e-04 pbeta0=-1.710825976e-11 agidl=2.635778408e-10 wagidl=-1.152507634e-15 bgidl=9.254056573e+08 lbgidl=8.270917627e+00 wbgidl=7.462837410e+03 pbgidl=-8.274690985e-4 cgidl=4.177955700e+02 lcgidl=-1.836079550e-05 wcgidl=-1.178493107e-02 pcgidl=1.836917206e-9 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.981765188e-01 lkt1=1.161947269e-08 wkt1=6.753731659e-06 pkt1=-1.162477373e-12 kt2=-3.805906314e-02 lkt2=-9.151132489e-10 wkt2=-5.637507627e-07 pkt2=9.155307419e-14 at=9.204209485e+04 lat=6.026373386e-04 wat=-1.142615893e-01 pat=-6.029122738e-8 ute=-2.110909566e-01 lute=8.271722411e-09 wute=4.449824834e-06 pute=-8.275496137e-13 ua1=1.959513039e-09 lua1=-2.581163689e-18 wua1=-1.243697535e-14 pua1=2.582341267e-22 ub1=-7.341682892e-19 lub1=8.199072311e-27 wub1=9.771284743e-24 pub1=-8.202812892e-31 uc1=-8.780780837e-11 luc1=1.993107584e-18 wuc1=1.549987650e-15 puc1=-1.994016880e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos lmin=2.0e-05 lmax=0.0001 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.102456397e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.153507141e-07 wvth0=-5.040651754e-08 pvth0=5.040090729e-12 k1=4.350633756e-01 lk1=1.508276488e-07 wk1=1.062792890e-08 pk1=-1.062674601e-12 k2=3.028188102e-02 lk2=-2.494815317e-07 wk2=-1.757948228e-08 pk2=1.757752569e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.323840640e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.996850373e-07 wvoff=2.111702525e-08 pvoff=-2.111467492e-12 nfactor='7.636495380e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.091700685e-05 wnfactor=7.692566545e-07 pnfactor=-7.691710363e-11 eta0=0.08 etab=-0.07 u0=1.618350503e-02 lu0=3.423211929e-07 wu0=2.412134198e-08 pu0=-2.411865728e-12 ua=-4.980122662e-10 lua=2.215036401e-14 wua=1.560804637e-15 pua=-1.560630920e-19 ub=2.018945184e-18 lub=3.248703844e-23 wub=2.289168712e-24 pub=-2.288913927e-28 uc=-7.885964217e-11 luc=1.188813844e-16 wuc=8.376865321e-18 puc=-8.375932976e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.749829144e+05 lvsat=2.501430123e+00 wvsat=1.762609289e-01 pvsat=-1.762413111e-5 a0=1.608197513e+00 la0=-1.066327438e-05 wa0=-7.513776341e-07 pa0=7.512940058e-11 ags=4.605314300e-01 lags=-7.864057630e-06 wags=-5.541334496e-07 pags=5.540717745e-11 a1=0.0 a2=8.739259507e-01 la2=1.260500183e-05 wa2=8.881996389e-07 pa2=-8.881007823e-11 b0=0.0 b1=0.0 keta=-3.644330552e-02 lketa=2.327163310e-06 wketa=1.639813812e-07 pketa=-1.639631301e-11 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.385060400e-01 lpclm=-6.300936432e-06 wpclm=-4.439895795e-07 ppclm=4.439401635e-11 pdiblc1=0.39 pdiblc2=1.445818285e-03 lpdiblc2=2.181538282e-07 wpdiblc2=1.537200502e-08 ppdiblc2=-1.537029412e-12 pdiblcb=-1.967595829e-03 lpdiblcb=1.871643453e-07 wpdiblcb=1.318836015e-08 ppdiblcb=-1.318689229e-12 drout=0.56 pscbe1=7.289941771e+08 lpscbe1=1.747900731e+03 wpscbe1=1.231641866e+02 ppscbe1=-1.231504784e-2 pscbe2=9.567980904e-09 lpscbe2=-6.298139368e-15 wpscbe2=-4.437924870e-16 ppscbe2=4.437430929e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=3.360966458e-10 lalpha0=-2.360703682e-14 walpha0=-1.663447722e-15 palpha0=1.663262580e-19 alpha1=3.713834012e-11 lalpha1=6.285466338e-15 walpha1=4.428994938e-16 palpha1=-4.428501991e-20 beta0=3.797941871e+00 lbeta0=9.943365472e-05 wbeta0=7.006499276e-06 pbeta0=-7.005719452e-10 agidl=3.216637424e-09 lagidl=-2.528236000e-13 wagidl=-1.781497799e-14 pagidl=1.781299518e-18 bgidl=1.341006471e+09 lbgidl=-1.865411064e+04 wbgidl=-1.314444421e+03 pbgidl=1.314298123e-1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.353864824e-01 lkt1=-6.302816058e-07 wkt1=-4.441220256e-08 pkt1=4.440725948e-12 kt2=-0.037961 at=0.0 ute=-3.322217128e-01 lute=3.155820000e-06 wute=2.223718982e-07 pute=-2.223471482e-11 ua1=2.2116e-9 ub1=-8.736257635e-19 lub1=8.002685548e-24 wub1=5.639017359e-25 pub1=-5.638389736e-29 uc1=1.1985e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.138243848e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' wvth0=2.017383375e-7 k1=4.426089572e-01 wk1=-4.253538653e-8 k2=1.780085875e-02 wk2=7.035708285e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.173914687e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' wvoff=-8.451513366e-8 nfactor='8.182649657e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=-3.078739937e-6 eta0=0.08 etab=-0.07 u0=3.330909506e-02 wu0=-9.653909194e-8 ua=6.101226114e-10 wua=-6.246694835e-15 ub=3.644201561e-18 wub=-9.161773375e-24 uc=-7.291226324e-11 wuc=-3.352611857e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.001240616e+05 wvsat=-7.054362909e-1 a0=1.074736923e+00 wa0=3.007184034e-6 ags=6.710960921e-02 wags=2.217767986e-6 a1=0.0 a2=1.504526972e+00 wa2=-3.554776789e-6 b0=0.0 b1=0.0 keta=7.997964934e-02 wketa=-6.562907508e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.767162027e-01 wpclm=1.776947189e-6 pdiblc1=0.39 pdiblc2=1.235958321e-02 wpdiblc2=-6.152225722e-8 pdiblcb=7.395832182e-03 wpdiblcb=-5.278281424e-8 drout=0.56 pscbe1=8.164378760e+08 wpscbe1=-4.929310625e+2 pscbe2=9.252898593e-09 wpscbe2=1.776158380e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-8.449124269e-10 walpha0=6.657495783e-15 alpha1=3.515866475e-10 walpha1=-1.772584419e-15 beta0=8.772392889e+00 wbeta0=-2.804160225e-5 agidl=-9.431581308e-09 wagidl=7.129959017e-14 bgidl=4.077815992e+08 wbgidl=5.260705265e+3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.669181100e-01 wkt1=1.777477268e-7 kt2=-0.037961 at=0.0 ute=-1.743428532e-01 wute=-8.899828683e-7 ua1=2.2116e-9 ub1=-4.732686873e-19 wub1=-2.256862888e-24 uc1=1.1985e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.161307916e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.842558420e-07 wvth0=2.821421361e-07 pvth0=-6.423354941e-13 k1=6.151870697e-01 lk1=-1.378704106e-06 wk1=-1.210094400e-06 pk1=9.327477176e-12 k2=-5.761121188e-02 lk2=6.024572286e-07 wk2=5.640866218e-07 pk2=-3.944341102e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.047521900e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.009735549e-07 wvoff=-2.541187408e-07 pvoff=1.354941169e-12 nfactor='8.922471357e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.910339387e-06 wnfactor=-6.339050955e-06 pnfactor=2.604620088e-11 eta0=0.08 etab=-0.07 u0=4.409550313e-02 lu0=-8.617121182e-08 wu0=-1.462604546e-07 pu0=3.972175026e-13 ua=1.689467794e-09 lua=-8.622748347e-15 wua=-1.146320274e-14 pua=4.167400354e-20 ub=4.242766131e-18 lub=-4.781854536e-24 wub=-1.157016041e-23 pub=1.924029091e-29 uc=-1.289764046e-10 luc=4.478891366e-16 wuc=3.105199470e-16 puc=-2.748539291e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.978419404e+05 lvsat=-7.806554309e-01 wvsat=-8.720088870e-01 pvsat=1.330726816e-6 a0=3.124989687e-01 la0=6.089419929e-06 wa0=6.251489093e-06 pa0=-2.591833136e-11 ags=-5.254099780e-01 lags=4.733561955e-06 wags=4.620952816e-06 pags=-1.919873119e-11 a1=0.0 a2=2.207093597e+00 la2=-5.612713438e-06 wa2=-7.099662412e-06 pa2=2.831963040e-11 b0=0.0 b1=0.0 keta=2.245044653e-01 lketa=-1.154589967e-06 wketa=-1.377977688e-06 pketa=5.765463121e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-9.839923918e-01 lpclm=6.449224529e-06 wpclm=3.548950023e-06 ppclm=-1.415630028e-11 pdiblc1=0.39 pdiblc2=2.354622109e-02 lpdiblc2=-8.936859575e-08 wpdiblc2=-1.182104019e-07 ppdiblc2=4.528742185e-13 pdiblcb=9.804416972e-03 lpdiblcb=-1.924187077e-08 wpdiblcb=-6.500789127e-08 ppdiblcb=9.766455109e-14 drout=0.56 pscbe1=6.416216750e+08 lpscbe1=1.396583904e+03 wpscbe1=3.626911329e+02 ppscbe1=-6.835454488e-3 pscbe2=9.812222954e-09 lpscbe2=-4.468369613e-15 wpscbe2=1.730604322e-15 ppscbe2=3.639254470e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-1.787195635e-09 lalpha0=7.527778052e-15 walpha0=1.329646708e-14 palpha0=-5.303787866e-20 alpha1=6.024732552e-10 lalpha1=-2.004300493e-15 walpha1=-3.540236621e-15 palpha1=1.412154365e-20 beta0=1.385922935e+01 lbeta0=-4.063807519e-05 wbeta0=-6.756341667e-05 pbeta0=3.157346375e-10 agidl=3.039339787e-06 lagidl=-2.435623812e-11 wagidl=-2.140612719e-11 pagidl=1.715803705e-16 bgidl=2.400996867e+09 lbgidl=-1.592353766e+04 wbgidl=-7.697605605e+03 pbgidl=1.035222610e-1 cgidl=300.0 egidl=6.277691851e-01 legidl=-4.216279410e-06 wegidl=-3.718462182e-06 pegidl=2.970631097e-11 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.390203810e-01 lkt1=-2.228713302e-07 wkt1=5.686108277e-08 pkt1=9.657476841e-13 kt2=-4.616153859e-02 lkt2=6.551303671e-08 wkt2=7.453494696e-08 pkt2=-5.954500017e-13 at=-4.616340251e+05 lat=3.687934214e+00 wat=1.408098974e+00 pat=-1.124911965e-5 ute=-2.299268933e+00 lute=1.697575821e-05 wute=1.406451037e-05 pute=-1.194695024e-10 ua1=-4.928623343e-09 lua1=5.704231605e-14 wua1=4.885433424e-14 pua1=-3.902909252e-19 ub1=4.325482046e-18 lub1=-3.833659577e-23 wub1=-3.484290359e-23 pub1=2.603256430e-28 uc1=-8.907706144e-11 luc1=1.669091133e-15 wuc1=1.352086981e-15 puc1=-1.080164712e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.116408964e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=5.159759037e-09 wvth0=9.292603865e-08 pvth0=1.124229204e-13 k1=1.423484992e-01 lk1=5.073874829e-07 wk1=1.567950669e-06 pk1=-1.753783457e-12 k2=1.499335278e-01 lk2=-2.254117573e-07 wk2=-6.363463596e-07 pk2=8.440300048e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.293770610e+00 ldsub=-2.926915574e-06 wdsub=-3.702329134e-06 pdsub=1.476810961e-11 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.562469675e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.044324184e-07 wvoff=-1.744421764e-07 pvoff=1.037121712e-12 nfactor='6.149705994e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=5.149861188e-06 wnfactor=1.116627186e-05 pnfactor=-4.378025612e-11 eta0=3.585049213e-01 leta0=-1.110919925e-06 weta0=-1.405230558e-06 peta0=5.605282015e-12 etab=-3.134728557e-01 letab=9.711815699e-07 wetab=1.228471997e-06 petab=-4.900215095e-12 u0=2.594602500e-02 lu0=-1.377530300e-08 wu0=-4.944853859e-08 pu0=1.104735514e-14 ua=-5.138352943e-10 lua=1.659412420e-16 wua=1.152263293e-15 pua=-8.647450472e-21 ub=3.707973304e-18 lub=-2.648635473e-24 wub=-9.976797850e-24 pub=1.288457481e-29 uc=7.129056065e-11 luc=-3.509497529e-16 wuc=-9.818053309e-16 puc=2.406378240e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.928848552e+05 lvsat=-3.619952623e-01 wvsat=-6.962348514e-01 pvsat=6.295870386e-7 a0=1.740018722e+00 la0=3.952292115e-07 wa0=6.870056538e-07 pa0=-3.722330298e-12 ags=5.840286448e-01 lags=3.081555154e-07 wags=-8.590439022e-07 pags=2.660263319e-12 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.730298644e-02 lketa=8.916942351e-08 wketa=2.410822573e-07 pketa=-6.927565222e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.735829217e-01 lpclm=1.432920088e-06 wpclm=2.697257863e-06 ppclm=-1.075901097e-11 pdiblc1=0.39 pdiblc2=1.962187643e-03 lpdiblc2=-3.272692266e-09 wpdiblc2=-8.815648409e-09 ppdiblc2=1.651276809e-14 pdiblcb=1.145869460e-02 lpdiblcb=-2.584056916e-08 wpdiblcb=-8.078046494e-08 ppdiblcb=1.605792971e-13 drout=0.56 pscbe1=1.181086351e+09 lpscbe1=-7.552705583e+02 wpscbe1=-2.684990378e+03 ppscbe1=5.321350861e-3 pscbe2=9.692068049e-09 lpscbe2=-3.989087317e-15 wpscbe2=-3.275750079e-15 ppscbe2=2.033362233e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=2.780816322e-03 lalpha0=-1.109231440e-08 walpha0=-1.959257995e-08 palpha0=7.815225438e-14 alpha1=-1.508771557e-10 lalpha1=1.000716360e-15 walpha1=1.767585607e-15 palpha1=-7.050669202e-21 beta0=6.776916852e+01 lbeta0=-2.556778142e-04 wbeta0=-4.538596138e-04 pbeta0=1.856619949e-9 agidl=-6.111699565e-06 lagidl=1.214606822e-11 wagidl=4.306250069e-11 pagidl=-8.557660520e-17 bgidl=-3.329181833e+09 lbgidl=6.933400255e+03 wbgidl=3.050177876e+04 pbgidl=-4.885011737e-2 cgidl=300.0 egidl=-9.555383702e-01 legidl=2.099328598e-06 wegidl=7.436924363e-06 pegidl=-1.479107576e-11 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.882472553e-01 lkt1=3.723752719e-07 wkt1=8.040359317e-07 pkt1=-2.014635656e-12 kt2=-2.943788167e-02 lkt2=-1.195456665e-09 wkt2=-5.339700739e-08 pkt2=-8.514606699e-14 at=7.379216042e+05 lat=-1.096937249e+00 wat=-2.147199903e+00 pat=2.932505380e-6 ute=4.316411536e+00 lute=-9.413331140e-06 wute=-3.343546404e-05 pute=7.000172055e-11 ua1=1.787229139e-08 lua1=-3.390756870e-14 wua1=-1.047961370e-13 pua1=2.226008302e-19 ub1=-1.147124632e-17 lub1=2.467450012e-23 wub1=7.168180679e-23 pub1=-1.645875785e-28 uc1=1.047266131e-09 luc1=-2.863634138e-15 wuc1=-4.947967883e-15 puc1=1.432845273e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.151608580e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=7.516721855e-08 wvth0=2.677413534e-07 pvth0=-2.352620146e-13 k1=3.426293699e-01 lk1=1.090548675e-07 wk1=1.422595963e-06 pk1=-1.464691844e-12 k2=4.309155025e-02 lk2=-1.291695333e-08 wk2=-3.964417812e-07 pk2=3.668909860e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.708461534e+00 ldsub=3.044133870e-06 wdsub=9.982070188e-06 pdsub=-1.244838167e-11 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.958003270e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.578809147e-08 wvoff=2.576265907e-07 pvoff=1.777931027e-13 nfactor='1.128424307e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.062065562e-06 wnfactor=-1.612127335e-05 pnfactor=1.049112392e-11 eta0=-6.146900923e-01 leta0=8.246384413e-07 weta0=2.806618621e-06 peta0=-2.771538461e-12 etab=-4.063511457e-01 letab=1.155904414e-06 wetab=2.862957363e-06 petab=-8.150994004e-12 u0=2.492582962e-02 lu0=-1.174626702e-08 wu0=-7.655926272e-08 pu0=6.496706104e-14 ua=1.764193197e-10 lua=-1.206885452e-15 wua=-8.093219902e-15 pua=9.740613691e-21 ub=2.635229046e-18 lub=-5.150866001e-25 wub=-2.792691989e-24 pub=-1.403677816e-30 uc=-1.277722590e-10 luc=4.496031725e-17 wuc=3.259101763e-16 puc=-1.944979013e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.273593820e+04 lvsat=3.607491425e-02 wvsat=-4.731944871e-01 pvsat=1.859887492e-7 a0=6.583297930e-01 la0=2.546567871e-06 wa0=7.730086770e-06 pa0=-1.773010304e-11 ags=-4.065775903e-01 lags=2.278342538e-06 wags=7.728853142e-06 pags=-1.441994747e-11 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=2.766171263e-02 lketa=-1.394804175e-07 wketa=-7.111568984e-07 pketa=1.201123367e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.689760276e-01 lpclm=4.987360150e-08 wpclm=-3.322450308e-06 ppclm=1.213406018e-12 pdiblc1=5.326869814e-01 lpdiblc1=-2.837858568e-07 wpdiblc1=-6.886815378e-07 ppdiblc1=1.369698050e-12 pdiblc2=2.046297715e-04 lpdiblc2=2.228618578e-10 wpdiblc2=-1.020410556e-09 ppdiblc2=1.009053386e-15 pdiblcb=-6.075014542e-02 lpdiblcb=1.177734265e-07 wpdiblcb=4.157835738e-07 ppdiblcb=-8.270220226e-13 drout=-9.238901618e-02 ldrout=1.297516943e-06 wdrout=2.580118768e-06 pdrout=-5.131520814e-12 pscbe1=8.026606526e+08 lpscbe1=-2.631039524e+00 wpscbe1=-1.874595240e+01 ppscbe1=1.853730995e-5 pscbe2=6.547310944e-09 lpscbe2=2.265425748e-15 wpscbe2=1.196539533e-14 ppscbe2=-9.979034533e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-5.526342102e-03 lalpha0=5.429543773e-09 walpha0=3.893651820e-08 palpha0=-3.825451305e-14 alpha1=3.522811000e-10 walpha1=-1.777477268e-15 beta0=-8.153451963e+01 lbeta0=4.126781201e-05 wbeta0=6.152475333e-04 pbeta0=-2.696951824e-10 agidl=-2.882044139e-09 lagidl=-3.575683908e-15 wagidl=1.983922098e-14 pagidl=2.965291472e-20 bgidl=-1.206890748e+08 lbgidl=5.521252629e+02 wbgidl=7.014341783e+03 pbgidl=-2.136658580e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.551411609e-01 lkt1=-9.124244614e-08 wkt1=-2.520107908e-07 pkt1=8.570398938e-14 kt2=-1.154294599e-02 lkt2=-3.678615740e-08 wkt2=-2.021935746e-07 pkt2=2.107909617e-13 at=1.326236721e+05 lat=1.069216493e-01 wat=-6.807401875e-01 pat=1.590764569e-8 ute=5.080731928e-01 lute=-1.839041260e-06 wute=3.913726864e-06 pute=-4.280964767e-12 ua1=2.914363291e-09 lua1=-4.158194237e-15 wua1=9.676223884e-15 pua1=-5.069814264e-21 ub1=6.859052361e-23 lub1=1.859546029e-24 wub1=-1.424483372e-23 pub1=6.309338986e-30 uc1=-6.961398448e-10 luc1=6.037737057e-16 wuc1=3.893070716e-15 puc1=-3.255223712e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.046727681e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.854635615e-08 wvth0=-2.842716136e-07 pvth0=3.106070481e-13 k1=4.367941770e-01 lk1=1.593811473e-08 wk1=-1.847848047e-07 pk1=1.247987759e-13 k2=4.316230198e-02 lk2=-1.298691759e-08 wk2=-4.659581481e-08 pk2=2.093880519e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.731635027e+00 ldsub=-3.576744154e-07 wdsub=-5.154823839e-06 pdsub=2.520038730e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.439872086e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.186247016e-08 wvoff=3.947914195e-07 pvoff=4.215491846e-14 nfactor='6.526113617e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.568940926e-07 wnfactor=-2.749870340e-06 pnfactor=-2.731455379e-12 eta0=5.200509789e-01 leta0=-2.974729618e-07 weta0=-6.992748246e-07 peta0=6.953343906e-13 etab=1.511287979e+00 letab=-7.403913865e-07 wetab=-1.065500945e-05 petab=5.216517842e-12 u0=1.283188478e-02 lu0=2.130722221e-10 wu0=8.999456157e-09 pu0=-1.963938929e-14 ua=-1.736210452e-09 lua=6.844567498e-16 wua=7.704838107e-15 pua=-5.881611933e-21 ub=3.124040065e-18 lub=-9.984571528e-25 wub=-9.132687820e-24 pub=4.865753860e-30 uc=-1.379956254e-10 luc=5.506989761e-17 wuc=1.835153721e-16 puc=-5.368795118e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.354245624e+05 lvsat=-1.050255855e-01 wvsat=-8.090486941e-01 pvsat=5.181048989e-7 a0=5.791699369e+00 la0=-2.529667301e-06 wa0=-2.338723892e-05 pa0=1.304088682e-11 ags=3.247094524e+00 lags=-1.334664206e-06 wags=-1.643481980e-05 pags=9.474783784e-12 a1=0.0 a2=1.883321980e-01 la2=6.048599394e-07 wa2=2.931891719e-06 pa2=-2.899259765e-12 b0=0.0 b1=0.0 keta=-1.978374128e-01 lketa=8.350890261e-08 wketa=1.021553884e-06 pketa=-5.123023442e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.098471692e-01 lpclm=5.038923557e-07 wpclm=3.434340253e-07 ppclm=-2.411677023e-12 pdiblc1=1.271271525e+00 lpdiblc1=-1.014149954e-06 wpdiblc1=-4.540081969e-06 ppdiblc1=5.178232394e-12 pdiblc2=2.136751842e-03 lpdiblc2=-1.687755694e-09 wpdiblc2=-1.441310473e-08 ppdiblc2=1.425268687e-14 pdiblcb=1.398423604e-01 lpdiblcb=-8.058648472e-08 wpdiblcb=-8.317322400e-07 ppdiblcb=4.066089402e-13 drout=8.712825320e-01 ldrout=3.445710587e-07 wdrout=-8.693426349e-07 pdrout=-1.720451917e-12 pscbe1=9.413387817e+08 lpscbe1=-1.397656810e+02 wpscbe1=-7.131420662e+02 ppscbe1=7.052047950e-4 pscbe2=8.935615814e-09 lpscbe2=-9.629728971e-17 wpscbe2=9.730156006e-16 ppscbe2=8.910000061e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-7.058038197e-05 lalpha0=3.450468022e-11 walpha0=4.972833965e-10 palpha0=-2.431069341e-16 alpha1=5.989464227e-10 lalpha1=-2.439199377e-16 walpha1=-3.515387893e-15 palpha1=1.718567679e-21 beta0=-8.738881919e+01 lbeta0=4.705695321e-05 wbeta0=6.760164052e-04 pbeta0=-3.297876966e-10 agidl=-1.365151909e-08 lagidl=7.073926786e-15 wagidl=9.896600536e-14 pagidl=-4.859318855e-20 bgidl=-2.886618402e+08 lbgidl=7.182284913e+02 wbgidl=9.677666015e+03 pbgidl=-4.770340014e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.077320673e-01 lkt1=-3.923687649e-08 wkt1=-3.105783279e-07 pkt1=1.436196698e-13 kt2=-6.831870466e-02 lkt2=1.935768709e-08 wkt2=4.885926778e-08 pkt2=-3.746766260e-14 at=4.632962301e+05 lat=-2.200705231e-01 wat=-1.499581909e+00 pat=8.256356592e-7 ute=-2.565694443e+00 lute=1.200515342e-06 wute=-8.215953660e-07 pute=4.016533266e-13 ua1=-5.201764567e-09 lua1=3.867601118e-15 wua1=9.982821821e-15 pua1=-5.372999766e-21 ub1=6.150217945e-18 lub1=-4.222152163e-24 wub1=-1.832412900e-23 pub1=1.034323171e-29 uc1=5.474096425e-11 luc1=-1.387498000e-16 wuc1=9.565556876e-16 puc1=-3.513920959e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.124905128e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=9.672252686e-09 wvth0=5.192623469e-07 pvth0=-8.221659921e-14 k1=2.357404101e-01 lk1=1.142272698e-07 wk1=-8.598265993e-08 pk1=7.649737133e-14 k2=9.900206785e-02 lk2=-4.028530393e-08 wk2=2.648302626e-08 pk2=-1.478724785e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.394750045e+00 ldsub=-1.929814546e-07 wdsub=-6.507213452e-07 pdsub=3.181181441e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.843516210e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.004824204e-07 wvoff=1.086841248e-06 pvoff=-2.961674811e-13 nfactor='7.496109875e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-8.310961629e-07 wnfactor=-1.127449939e-05 pnfactor=1.435980024e-12 eta0=-6.411277589e-01 leta0=2.701924878e-07 weta0=1.413919628e-06 peta0=-3.377429816e-13 etab=-5.674954363e-03 letab=1.206282599e-09 wetab=3.041347972e-08 petab=-7.264867901e-15 u0=2.091693257e-02 lu0=-3.739465095e-09 wu0=-6.138745316e-08 pu0=1.477065907e-14 ua=1.245578941e-09 lua=-7.732506304e-16 wua=-9.535092306e-15 pua=2.546472848e-21 ub=2.762732061e-19 lub=3.937306315e-25 wub=2.510336035e-24 pub=-8.261712118e-31 uc=-8.230069429e-11 luc=2.784231663e-17 wuc=3.745930698e-16 puc=-1.471001053e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.929130848e+04 lvsat=2.927476224e-02 wvsat=5.803532862e-01 pvsat=-1.611320472e-7 a0=3.687733935e-01 la0=1.214385206e-07 wa0=7.071224328e-06 pa0=-1.849342110e-12 ags=-2.019838439e+00 lags=1.240181312e-06 wags=1.158989026e-05 pags=-4.225656222e-12 a1=0.0 a2=2.023335604e+00 la2=-2.922181757e-07 wa2=-5.863783439e-06 pa2=1.400681950e-12 b0=0.0 b1=0.0 keta=-2.775409284e-04 lketa=-1.307219194e-08 wketa=1.671825008e-07 pketa=-9.462580599e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.119052267e+00 lpclm=-2.827997406e-07 wpclm=-7.541388585e-06 ppclm=1.442976206e-12 pdiblc1=-2.057828753e+00 lpdiblc1=6.133472987e-07 wpdiblc1=1.274411926e-05 ppdiblc1=-3.271495060e-12 pdiblc2=-1.052193208e-02 lpdiblc2=4.500695113e-09 wpdiblc2=2.780959603e-08 ppdiblc2=-6.388724848e-15 pdiblcb=-0.025 drout=2.260665214e+00 ldrout=-3.346564528e-07 wdrout=-6.578929859e-06 pdrout=1.070793990e-12 pscbe1=5.173224367e+08 lpscbe1=6.752318955e+01 wpscbe1=1.426284132e+03 ppscbe1=-3.406964907e-4 pscbe2=1.613274885e-08 lpscbe2=-3.614759719e-15 wpscbe2=5.466712571e-15 ppscbe2=-1.305833632e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-5.268145045e-08 lalpha0=2.580326768e-14 walpha0=2.663152476e-13 palpha0=-1.301935351e-19 alpha1=4.365975454e-10 lalpha1=-1.645524420e-16 walpha1=-1.698343980e-15 palpha1=8.302694217e-22 beta0=-1.744304970e+01 lbeta0=1.286256489e-05 wbeta0=1.357789499e-04 pbeta0=-6.568181191e-11 agidl=-3.000597701e-10 lagidl=5.467988687e-16 wagidl=4.343938651e-15 pagidl=-2.335298802e-21 bgidl=1.015572358e+09 lbgidl=8.062751900e+01 wbgidl=5.891334639e+02 pbgidl=-3.272291055e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.325448675e-01 lkt1=-2.710664286e-08 wkt1=-3.636361277e-07 pkt1=1.695580364e-13 kt2=-2.386568597e-02 lkt2=-2.374060162e-09 wkt2=-2.358096856e-08 pkt2=-2.053804258e-15 at=-3.680751891e+04 lat=2.441519666e-02 wat=5.055652706e-01 pat=-1.546206427e-7 ute=-1.118874046e-01 lute=9.226954631e-10 wute=-3.906191155e-07 pute=1.909619670e-13 ua1=4.214192790e-09 lua1=-7.355779551e-16 wua1=-2.430299690e-15 pua1=6.954029476e-22 ub1=-4.504795523e-18 lub1=9.867642713e-25 wub1=8.025112197e-24 pub1=-2.538121832e-30 uc1=-3.249743350e-10 luc1=4.688161836e-17 wuc1=9.759192973e-17 puc1=6.852951647e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.025480288e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.344218766e-08 wvth0=4.540308671e-07 pvth0=-6.663475565e-14 k1=-4.824469119e-01 lk1=2.857806754e-07 wk1=4.636705560e-06 pk1=-1.051611164e-12 k2=3.316496711e-01 lk2=-9.585783692e-08 wk2=-1.452378614e-06 pk2=3.384684322e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.287085407e+00 ldsub=-6.450036024e-07 wdsub=-1.632919047e-05 pdsub=4.063234064e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.799512326e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.883299661e-09 wvoff=-5.006072347e-08 pvoff=-2.459570722e-14 nfactor='5.143933348e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.692317559e-07 wnfactor=-1.472090504e-05 pnfactor=2.259222941e-12 eta0=0.49 etab=-6.249997450e-04 letab=-6.090131524e-17 wetab=-1.286411089e-15 petab=3.072850160e-22 u0=2.030169749e-02 lu0=-3.592503891e-09 wu0=-7.451192946e-08 pu0=1.790570272e-14 ua=1.888973283e-09 lua=-9.269382369e-16 wua=-2.064889989e-14 pua=5.201228065e-21 ub=-3.001704319e-19 lub=5.314257234e-25 wub=1.346828750e-23 pub=-3.443697078e-30 uc=6.421360169e-11 luc=-7.155553250e-18 wuc=-2.659910428e-16 puc=5.916221718e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.789257656e+05 lvsat=-2.285075025e-02 wvsat=-7.984992117e-01 pvsat=1.682344489e-7 a0=3.322190226e+00 la0=-5.840441581e-07 wa0=-1.488909283e-05 pa0=3.396318850e-12 ags=7.808785771e+00 lags=-1.107582153e-06 wags=-2.081684479e-05 pags=3.515340579e-12 a1=0.0 a2=3.954555545e-02 la2=1.816497532e-07 wa2=6.639653440e-06 pa2=-1.586014017e-12 b0=0.0 b1=0.0 keta=3.147414154e-01 lketa=-8.832077004e-08 wketa=-2.821847028e-06 pketa=6.193636776e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.187796882e+00 lpclm=-6.035076660e-08 wpclm=-2.958277732e-06 ppclm=3.482085171e-13 pdiblc1=8.626234743e-01 lpdiblc1=-8.426112488e-08 wpdiblc1=-3.993892463e-06 ppdiblc1=7.267138002e-13 pdiblc2=5.604675091e-03 lpdiblc2=6.485324593e-10 wpdiblc2=8.874469673e-09 ppdiblc2=-1.865691216e-15 pdiblcb=7.680222456e-01 lpdiblcb=-1.894292238e-07 wpdiblcb=-3.031142565e-06 ppdiblcb=7.240490246e-13 drout=5.179002047e-01 ldrout=8.163782487e-08 wdrout=-7.802466472e-08 pdrout=-4.820772341e-13 pscbe1=7.987271780e+08 lpscbe1=3.040389852e-01 wpscbe1=1.070594185e+01 ppscbe1=-2.557328329e-6 pscbe2=-5.473616084e-08 lpscbe2=1.331369674e-14 wpscbe2=2.519228739e-13 ppscbe2=-6.017681689e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=6.612550594e-08 lalpha0=-2.576149992e-15 walpha0=-3.331397454e-13 palpha0=1.299827908e-20 alpha1=-2.522811000e-10 walpha1=1.777477268e-15 beta0=4.221536133e+01 lbeta0=-1.388039759e-06 wbeta0=-1.722413283e-04 pbeta0=7.894991965e-12 agidl=6.546237020e-09 lagidl=-1.088576046e-15 wagidl=-1.853803110e-14 pagidl=3.130517311e-21 bgidl=-8.366471076e+08 lbgidl=5.230671827e+02 wbgidl=1.201349619e+04 pbgidl=-3.056166629e-3 cgidl=2.432791151e+03 lcgidl=-5.094598222e-04 wcgidl=-1.076125795e-02 pcgidl=2.570541687e-9 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-8.646056734e-01 lkt1=7.609972184e-08 wkt1=3.452081466e-07 pkt1=2.364046054e-16 kt2=1.271108929e-02 lkt2=-1.111115447e-08 wkt2=-1.098084317e-07 pkt2=1.854334986e-14 at=1.130772970e+05 lat=-1.138778932e-02 wat=-2.692591021e-01 pat=3.046165526e-8 ute=-1.407145244e+00 lute=3.103209356e-07 wute=1.154956856e-05 pute=-2.661190664e-12 ua1=2.961418227e-09 lua1=-4.363276953e-16 wua1=1.641103723e-15 pua1=-2.771331857e-22 ub1=-1.445563025e-18 lub1=2.560054044e-25 wub1=-8.873761167e-24 pub1=1.498512048e-30 uc1=-4.166419301e-10 luc1=6.877825681e-17 wuc1=1.312018582e-15 puc1=-2.215605779e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.022794758e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.546521643e-08 wvth0=-2.004391083e-07 pvth0=4.830351422e-14 k1=2.065713039e+00 lk1=-1.590765159e-07 wk1=-1.121392378e-05 pk1=1.788680505e-12 k2=-1.131625526e-01 lk2=-2.283051622e-08 wk2=2.137140567e-06 pk2=-2.946421674e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-5.065081894e+00 ldsub=8.424817669e-07 wdsub=4.902949247e-05 pdsub=-7.675941999e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.811061490e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.307589246e-08 wvoff=-1.054575633e-06 pvoff=1.596374499e-13 nfactor='1.229956199e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.626351784e-06 wnfactor=-2.058434267e-05 pnfactor=3.576494156e-12 eta0=1.891873008e+00 leta0=-2.605661360e-07 weta0=6.742604475e-09 peta0=-1.253247894e-15 etab=3.055636466e-01 letab=-5.691128375e-08 wetab=-8.676670805e-07 petab=1.612732803e-13 u0=-3.532497796e-02 lu0=6.385171948e-09 wu0=2.495363411e-07 pu0=-4.052259739e-14 ua=-1.465795725e-08 lua=2.055325654e-15 wua=7.970326381e-14 pua=-1.292762537e-20 ub=1.121124418e-17 lub=-1.554702733e-24 wub=-5.765139062e-23 pub=9.428643424e-30 uc=2.753551710e-10 luc=-4.712078022e-17 wuc=-1.868166604e-15 puc=3.043081744e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.545274462e+04 lvsat=1.469541776e-02 wvsat=1.315064650e+00 pvsat=-2.076776465e-7 a0=-7.273413919e-01 la0=1.098470525e-07 wa0=9.823905579e-06 pa0=-8.551816199e-13 ags=1.25 a1=0.0 a2=2.924370978e+00 la2=-3.362662212e-07 wa2=-1.766774448e-05 pa2=2.772339345e-12 b0=-3.857065301e-23 lb0=7.169127274e-30 wb0=1.946129354e-28 pb0=-3.617270630e-35 b1=0.0 keta=-1.000116229e+00 lketa=1.471806431e-07 wketa=3.989826405e-06 pketa=-5.843712461e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.867697356e+00 lpclm=-1.927993284e-07 wpclm=-5.446429493e-06 ppclm=8.457351416e-13 pdiblc1=9.676613367e-01 lpdiblc1=-1.122670085e-07 wpdiblc1=4.436304055e-06 ppdiblc1=-7.670491633e-13 pdiblc2=3.218940421e-02 lpdiblc2=-4.227483929e-09 wpdiblc2=3.086863098e-08 ppdiblc2=-6.141563533e-15 pdiblcb=-2.420745796e+00 lpdiblcb=3.841974125e-07 wpdiblcb=1.557684790e-05 ppdiblcb=-2.661728760e-12 drout=1.008278222e+00 ldrout=-1.290326457e-09 wdrout=-1.817033286e-05 pdrout=2.832209783e-12 pscbe1=8.032688971e+08 lpscbe1=-5.095229859e-01 wpscbe1=-2.749529989e+01 ppscbe1=4.285692394e-6 pscbe2=9.832662827e-08 lpscbe2=-1.379580529e-14 wpscbe2=-6.358906359e-13 ppscbe2=9.878313094e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=2.133641271e-07 lalpha0=-3.020273135e-14 walpha0=-1.076050171e-12 palpha0=1.523915657e-19 alpha1=-2.522811000e-10 walpha1=1.777477268e-15 beta0=6.333469369e+01 lbeta0=-5.453222852e-06 wbeta0=-2.466382006e-04 pbeta0=2.251792078e-11 agidl=1.0e-10 bgidl=4.621900562e+09 lbgidl=-4.388563421e+02 wbgidl=-1.858126842e+04 pbgidl=2.322820559e-3 cgidl=-5.177494006e+03 lcgidl=8.537769907e-04 wcgidl=2.763736426e-02 pcgidl=-4.307835967e-9 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=3.516767462e-01 lkt1=-1.423097969e-07 wkt1=7.659867988e-07 pkt1=-7.794992482e-14 kt2=-7.634695936e-01 lkt2=1.320389985e-07 wkt2=4.547217630e-06 pkt2=-8.451913409e-13 at=4.123296582e+05 lat=-6.815622480e-02 wat=-2.370886692e+00 pat=4.241577244e-7 ute=5.016015031e+00 lute=-8.523121187e-07 wute=-3.237838811e-05 pute=5.235798830e-12 ua1=-2.752956097e-09 lua1=5.818783204e-16 wua1=2.076530087e-14 pua1=-3.859646472e-21 ub1=4.684208350e-18 lub1=-8.575633536e-25 wub1=-2.840454891e-23 pub1=5.279553506e-30 uc1=4.806005855e-10 luc1=-9.106836066e-17 wuc1=-2.454803035e-15 puc1=4.562742401e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos lmin=2.0e-05 lmax=0.0001 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108794785e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-8.158245220e-08 wvth0=-1.842540719e-08 pvth0=1.842335644e-12 k1=4.568416918e-01 lk1=-2.026761573e-06 wk1=-9.925722216e-08 pk1=9.924617483e-12 k2=1.854189619e-02 lk2=9.243862853e-07 wk2=4.165604346e-08 pk2=-4.165140714e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.341091104e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.721704830e-07 wvoff=2.982095759e-08 pvoff=-2.981763851e-12 nfactor='7.958631595e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.129302935e-05 wnfactor=-8.561209224e-07 pnfactor=8.560256362e-11 eta0=0.08 etab=-0.07 u0=2.053201286e-02 lu0=-9.248119196e-08 wu0=2.180415171e-09 pu0=-2.180172491e-13 ua=-1.818148443e-10 lua=-9.465858904e-15 wua=-3.460803100e-17 pua=3.460417912e-21 ub=2.410868435e-18 lub=-6.700924611e-24 wub=3.116721315e-25 pub=-3.116374424e-29 uc=-8.847927211e-11 luc=1.080737311e-15 wuc=5.691388173e-17 puc=-5.690754722e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.099163535e+05 lvsat=-9.915249786e-1 a0=1.438607171e+00 la0=6.293872356e-06 wa0=1.043111304e-07 pa0=-1.042995206e-11 ags=3.399822733e-01 lags=4.189516329e-06 wags=5.411202764e-08 pags=-5.410600497e-12 a1=0.0 a2=1.049959676e+00 la2=-4.996411477e-6 b0=0.0 b1=0.0 keta=3.230853340e-03 lketa=-1.639811003e-06 wketa=-3.619942751e-08 pketa=3.619539852e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.635223146e-03 lpclm=6.884677536e-06 wpclm=2.213807154e-07 ppclm=-2.213560757e-11 pdiblc1=0.39 pdiblc2=4.538308903e-03 lpdiblc2=-9.106081414e-08 wpdiblc2=-2.315336763e-10 ppdiblc2=2.315079066e-14 pdiblcb=1.230263679e-03 lpdiblcb=-1.325860133e-07 wpdiblcb=-2.946830134e-09 ppdiblcb=2.946502152e-13 drout=0.56 pscbe1=7.806156748e+08 lpscbe1=-3.413674501e+03 wpscbe1=-1.372983783e+02 ppscbe1=1.372830970e-2 pscbe2=9.387039523e-09 lpscbe2=1.179398485e-14 wpscbe2=4.691693253e-16 ppscbe2=-4.691171067e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-1.360966458e-10 lalpha0=2.360703682e-14 walpha0=7.190611385e-16 palpha0=-7.189811070e-20 alpha1=1.628616599e-10 lalpha1=-6.285466338e-15 walpha1=-1.914528543e-16 palpha1=1.914315456e-20 beta0=5.104848607e+00 lbeta0=-3.124247305e-05 wbeta0=4.123418947e-07 pbeta0=-4.122960010e-11 agidl=-2.007477886e-09 lagidl=2.695297866e-13 wagidl=8.543933152e-15 pagidl=-8.542982212e-19 bgidl=9.091179662e+08 lbgidl=2.452993290e+04 wbgidl=8.647017195e+02 pbgidl=-8.646054782e-2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.532633165e-01 lkt1=1.157202834e-06 wkt1=4.578754482e-08 pkt1=-4.578244866e-12 kt2=-0.037961 at=0.0 ute=-2.801439377e-01 lute=-2.051377888e-06 wute=-4.039286973e-08 pute=4.038837400e-12 ua1=2.320991131e-09 lua1=-1.093789553e-14 wua1=-5.519462950e-16 pua1=5.518848634e-20 ub1=-1.051129558e-18 lub1=2.575108939e-23 wub1=1.459518787e-24 pub1=-1.459356343e-28 uc1=2.362916267e-10 luc1=-1.164286668e-14 wuc1=-5.875204336e-16 puc1=5.874550426e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.112876179e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' wvth0=7.374266654e-8 k1=3.554471871e-01 wk1=3.972499582e-7 k2=6.478694583e-02 wk2=-1.667169518e-7 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.104874408e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' wvoff=-1.193502488e-7 nfactor='6.893387320e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=3.426390476e-6 eta0=0.08 etab=-0.07 u0=1.590537854e-02 wu0=-8.726516991e-9 ua=-6.553713237e-10 wua=1.385092044e-16 ub=2.075635647e-18 wub=-1.247382695e-24 uc=-3.441231829e-11 wuc=-2.277822878e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160312.5 a0=1.753476013e+00 wa0=-4.174768475e-7 ags=5.495747279e-01 wags=-2.165686310e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-7.880534994e-02 wketa=1.448783348e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=3.510607727e-01 wpclm=-8.860159295e-7 pdiblc1=0.39 pdiblc2=-1.726698156e-05 wpdiblc2=9.266503862e-10 pdiblcb=-5.402728247e-03 wpdiblcb=1.179388383e-8 drout=0.56 pscbe1=6.098369114e+08 wpscbe1=5.494993096e+2 pscbe2=9.977067116e-09 wpscbe2=-1.877722254e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.044912427e-09 walpha0=-2.877846075e-15 alpha1=-1.515866475e-10 walpha1=7.662378286e-16 beta0=3.541855149e+00 wbeta0=-1.650285963e-6 agidl=1.147651529e-08 wagidl=-3.419476199e-14 bgidl=2.136297537e+09 wbgidl=-3.460732776e+3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.953709577e-01 wkt1=-1.832521591e-7 kt2=-0.037961 at=0.0 ute=-3.827699434e-01 wute=1.616614435e-7 ua1=1.773791837e-09 wua1=2.209014496e-15 ub1=2.371418346e-19 wub1=-5.841325846e-24 uc1=-3.461758503e-10 wuc1=2.351390283e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.122911590e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=8.017159459e-08 wvth0=8.840878645e-08 pvth0=-1.171657253e-13 k1=2.581902401e-01 lk1=7.769731063e-07 wk1=5.911766575e-07 pk1=-1.549255190e-12 k2=1.025307909e-01 lk2=-3.015306720e-07 wk2=-2.439293908e-07 pk2=6.168401374e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.286901560e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.454191253e-07 wvoff=-1.333368126e-07 pvoff=1.117368407e-13 nfactor='6.585697314e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.458095456e-06 wnfactor=5.451427567e-06 pnfactor=-1.617775807e-11 eta0=0.08 etab=-0.07 u0=1.359700336e-02 lu0=1.844130926e-08 wu0=7.623446800e-09 pu0=-1.306177352e-13 ua=-1.284830365e-09 lua=5.028666453e-15 wua=3.543981481e-15 pua=-2.720587530e-20 ub=2.417371494e-18 lub=-2.730083250e-24 wub=-2.359909068e-24 pub=8.887828571e-30 uc=4.661972086e-11 luc=-6.473544266e-16 wuc=-5.754717266e-16 puc=2.777645727e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.307415459e+05 lvsat=-5.626484918e-01 wvsat=-2.888346007e-02 pvsat=2.307462077e-7 a0=1.365375936e+00 la0=3.100481058e-06 wa0=9.390699015e-07 pa0=-1.083727563e-11 ags=2.907865540e-01 lags=2.067425079e-06 wags=5.027336373e-07 pags=-5.746412312e-12 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-6.559908778e-02 lketa=-1.055031116e-07 wketa=8.577518185e-08 pketa=4.721674059e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=7.009301966e-02 lpclm=2.244614854e-06 wpclm=-1.769566520e-06 ppclm=7.058570803e-12 pdiblc1=0.39 pdiblc2=-2.488876802e-04 lpdiblc2=1.850387651e-09 wpdiblc2=1.850722368e-09 ppdiblc2=-7.382290930e-15 pdiblcb=-7.090168188e-03 lpdiblcb=1.348073832e-08 wpdiblcb=2.023579930e-08 ppdiblcb=-6.744136523e-14 drout=0.56 pscbe1=6.114112903e+08 lpscbe1=-1.257750809e+01 wpscbe1=5.151213146e+02 ppscbe1=2.746413327e-4 pscbe2=1.168138527e-08 lpscbe2=-1.361557616e-14 wpscbe2=-7.700482174e-15 ppscbe2=4.651727205e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.987195635e-09 lalpha0=-7.527778052e-15 walpha0=-5.747684544e-15 palpha0=2.292676645e-20 alpha1=-4.024732552e-10 lalpha1=2.004300493e-15 walpha1=1.530343600e-15 palpha1=-6.104341677e-21 beta0=2.220999188e+00 lbeta0=1.055214657e-05 wbeta0=-8.841306526e-06 pbeta0=5.744812845e-11 agidl=-3.034768146e-06 lagidl=2.433605259e-11 wagidl=9.241525426e-12 pagidl=-7.410252274e-17 bgidl=9.867718769e+08 lbgidl=9.183411057e+03 wbgidl=-5.619608822e+02 pbgidl=-2.315791182e-2 cgidl=300.0 egidl=-4.277691851e-01 legidl=4.216279410e-06 wegidl=1.607385441e-06 pegidl=-1.284119333e-11 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.022916677e-01 lkt1=-7.435983468e-07 wkt1=-6.330203209e-07 pkt1=3.593139375e-12 kt2=-3.138933668e-02 lkt2=-5.250016399e-8 at=-1.881185878e+05 lat=1.502854942e+00 wat=2.804346631e-02 pat=-2.240356067e-7 ute=9.853518131e-01 lute=-1.092974686e-05 wute=-2.508444332e-06 pute=2.133112793e-11 ua1=3.879498199e-09 lua1=-1.682221438e-14 wua1=4.411882410e-15 pua1=-1.759842539e-20 ub1=-7.594419955e-20 lub1=2.501203626e-24 wub1=-1.263497049e-23 pub1=5.427354390e-29 uc1=-7.518597356e-10 luc1=3.240955820e-15 wuc1=4.696237823e-15 puc1=-1.873268216e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108410888e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.233017981e-08 wvth0=5.257076892e-08 pvth0=2.578746763e-14 k1=2.328244978e-01 lk1=8.781537546e-07 wk1=1.111442980e-06 pk1=-3.624529915e-12 k2=1.053904391e-01 lk2=-3.129374366e-07 wk2=-4.115987710e-07 pk2=1.285651498e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.897211863e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.888639712e-07 wvoff=-5.543921648e-09 pvoff=-3.980123885e-13 nfactor='8.273863182e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.275778731e-06 wnfactor=4.485776171e-07 pnfactor=3.777960013e-12 eta0=0.08 etab=-0.07 u0=2.832189895e-02 lu0=-4.029438503e-08 wu0=-6.143630048e-08 pu0=1.448526189e-13 ua=1.816042345e-09 lua=-7.340311674e-15 wua=-1.060341858e-14 pua=2.922626438e-20 ub=1.171029543e-18 lub=2.241412768e-24 wub=2.823661404e-24 pub=-1.178876018e-29 uc=-2.090983595e-10 luc=3.726717528e-16 wuc=4.329311734e-16 puc=-1.244742349e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.704228994e+05 lvsat=-3.220452523e-01 wvsat=-7.833811313e-02 pvsat=4.280143896e-7 a0=1.741545138e+00 la0=1.599991014e-06 wa0=6.793039346e-07 pa0=-9.801102954e-12 ags=5.764744137e-02 lags=2.997386691e-06 wags=1.796876678e-06 pags=-1.090858066e-11 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-3.699411678e-02 lketa=-2.196046222e-07 wketa=-1.275728226e-08 pketa=8.652005960e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.170973158e-01 lpclm=6.268582688e-08 wpclm=9.640140789e-07 ppclm=-3.845326839e-12 pdiblc1=0.39 pdiblc2=0.000215 pdiblcb=-4.139009881e-02 lpdiblcb=1.502987026e-07 wpdiblcb=1.858745697e-07 ppdiblcb=-7.281528875e-13 drout=0.56 pscbe1=4.189136490e+08 lpscbe1=7.552705583e+02 wpscbe1=1.160644974e+03 ppscbe1=-2.300268628e-3 pscbe2=-2.646401887e-09 lpscbe2=4.353610419e-14 wpscbe2=5.897950528e-14 ppscbe2=-2.194605295e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-2.780816122e-03 lalpha0=1.109231440e-08 walpha0=8.469315062e-09 palpha0=-3.378299677e-14 alpha1=3.508771557e-10 lalpha1=-1.000716360e-15 walpha1=-7.640769846e-16 palpha1=3.047803762e-21 beta0=-6.443688909e+01 lbeta0=2.764417974e-04 wbeta0=2.132021790e-04 pbeta0=-8.282544696e-10 agidl=6.111806933e-06 lagidl=-1.214844635e-11 wagidl=-1.861269262e-11 pagidl=3.700433199e-17 bgidl=5.111398910e+09 lbgidl=-7.269189978e+03 wbgidl=-1.208620113e+04 pbgidl=2.281078437e-2 cgidl=300.0 egidl=1.155538370e+00 legidl=-2.099328598e-06 wegidl=-3.214770882e-06 pegidl=6.393761365e-12 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.589575541e-01 lkt1=2.802085073e-07 wkt1=6.562511708e-07 pkt1=-1.549597000e-12 kt2=-3.978791304e-02 lkt2=-1.899933468e-08 wkt2=-1.174661393e-09 pkt2=4.685571591e-15 at=3.698768720e+05 lat=-7.229164073e-01 wat=-2.901853053e-01 pat=1.045337593e-6 ute=-3.330248395e+00 lute=6.284621347e-06 wute=5.146691534e-06 pute=-9.204213873e-12 ua1=-2.323147812e-09 lua1=7.919334216e-15 wua1=-2.897584698e-15 pua1=1.155808868e-20 ub1=2.073574380e-18 lub1=-6.072946550e-24 wub1=3.339761462e-24 pub1=-9.447585148e-30 uc1=2.772151415e-11 luc1=1.313075607e-16 wuc1=1.962688676e-16 puc1=-7.828909981e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.110269132e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.602598639e-08 wvth0=5.915812766e-08 pvth0=1.268606744e-14 k1=9.173808884e-01 lk1=-4.833399140e-07 wk1=-1.477382943e-06 pk1=1.524308298e-12 k2=-1.328242626e-01 lk2=1.608406371e-07 wk2=4.911629141e-07 pk2=-5.098241348e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.447643867e-02 ldsub=9.457545454e-07 wdsub=9.355829091e-07 pdsub=-1.860752781e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.028908370e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.728269429e-08 wvoff=-2.111595762e-07 pvoff=1.093041847e-14 nfactor='7.471656886e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.680294696e-06 wnfactor=3.115595359e-06 pnfactor=-1.526391564e-12 eta0=-5.995440838e-02 leta0=2.783511242e-07 weta0=7.632050099e-09 peta0=-1.517915548e-14 etab=-6.357158270e-01 letab=1.125135237e-06 wetab=4.020244845e-06 petab=-7.995744365e-12 u0=3.902060463e-03 lu0=8.273499145e-09 wu0=2.951872949e-08 pu0=-3.604511156e-14 ua=-3.309524365e-09 lua=2.853774189e-15 wua=9.495534245e-15 pua=-1.074793993e-20 ub=3.498445948e-18 lub=-2.387515897e-24 wub=-7.148158180e-24 pub=8.043892638e-30 uc=2.554573859e-11 luc=-9.400485470e-17 wuc=-4.476744853e-16 puc=5.066678276e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.413607529e+04 lvsat=1.444620556e-01 wvsat=3.183223954e-01 pvsat=-3.608917959e-7 a0=3.851883310e+00 la0=-2.597197266e-06 wa0=-8.383377113e-06 pa0=8.223391501e-12 ags=2.632588530e+00 lags=-2.123836391e-06 wags=-7.605630295e-06 pags=7.791783379e-12 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-2.817890151e-01 lketa=2.672606071e-07 wketa=8.502145011e-07 pketa=-8.511380948e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=7.207572630e-01 lpclm=-1.434803323e-07 wpclm=-2.070032248e-06 ppclm=2.188996880e-12 pdiblc1=3.769956971e-01 lpdiblc1=2.586386786e-08 wpdiblc1=9.687783153e-08 ppdiblc1=-1.926774128e-13 pdiblc2=2.392950000e-06 lpdiblc2=4.228477835e-10 pdiblcb=9.270092676e-02 lpdiblcb=-1.163909154e-07 wpdiblcb=-3.584725320e-07 ppdiblcb=3.544827327e-13 drout=8.523031487e-01 ldrout=-5.813529634e-07 wdrout=-2.186440802e-06 pdrout=4.348546518e-12 pscbe1=7.973393474e+08 lpscbe1=2.631039524e+00 wpscbe1=8.103342053e+00 ppscbe1=-8.013151856e-6 pscbe2=2.928315775e-08 lpscbe2=-1.996763908e-14 wpscbe2=-1.027510935e-13 ppscbe2=1.022006065e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=5.526342302e-03 lalpha0=-5.429543773e-09 walpha0=-1.683114939e-08 palpha0=1.653633796e-14 alpha1=-1.522811000e-10 walpha1=7.683528683e-16 beta0=9.158106374e+01 lbeta0=-3.385762846e-05 wbeta0=-2.582282627e-04 pbeta0=1.093593929e-10 agidl=1.667226227e-09 lagidl=3.827209458e-15 wagidl=-3.114677670e-15 pagidl=-7.699286911e-21 bgidl=1.270113134e+09 lbgidl=3.706280642e+02 wbgidl=-3.120438703e+00 pbgidl=-1.220892321e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.451299616e-01 lkt1=-1.450667767e-07 wkt1=-3.025235182e-07 pkt1=3.572812157e-13 kt2=-3.823071454e-02 lkt2=-2.209640007e-08 wkt2=-6.753718248e-08 pkt2=1.366719989e-13 at=-1.046632834e+05 lat=2.208822715e-01 wat=5.165200953e-01 pat=-5.590945767e-7 ute=3.238636071e+00 lute=-6.780035903e-06 wute=-9.863661269e-06 pute=2.064942651e-11 ua1=7.889564179e-09 lua1=-1.239242228e-14 wua1=-1.542675917e-14 pua1=3.647698791e-20 ub1=-4.796816849e-18 lub1=7.591368453e-24 wub1=9.958436984e-24 pub1=-2.261127033e-29 uc1=-4.245343738e-11 luc1=2.708764165e-16 wuc1=5.948161973e-16 puc1=-1.575549826e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.131892253e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.740844205e-08 wvth0=1.454366276e-07 pvth0=-7.263215276e-14 k1=5.026836058e-01 lk1=-7.325821210e-08 wk1=-5.172379558e-07 pk1=5.748497248e-13 k2=-7.579439947e-03 lk2=3.698978931e-08 wk2=2.094278346e-07 pk2=-2.312247666e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.080841523e+00 ldsub=-3.952099518e-08 wdsub=-1.871165818e-06 pdsub=9.147568336e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.114075640e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.570463012e-08 wvoff=-2.741553524e-07 pvoff=7.322505162e-14 nfactor='6.093805212e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.317778510e-06 wnfactor=-5.686055387e-07 pnfactor=2.116804178e-12 eta0=4.168013260e-01 leta0=-1.930983189e-07 weta0=-1.783161045e-07 peta0=1.686993961e-13 etab=9.925540395e-01 letab=-4.850119860e-07 wetab=-8.037674077e-06 petab=3.927969920e-12 u0=1.906757575e-02 lu0=-6.723223960e-09 wu0=-2.246348342e-08 pu0=1.535853932e-14 ua=3.717612460e-10 lua=-7.865387138e-16 wua=-2.931190266e-15 pua=1.540475141e-21 ub=1.347668433e-18 lub=-2.606765365e-25 wub=-1.697880345e-25 pub=1.143191751e-30 uc=-1.585804685e-10 luc=8.807202769e-17 wuc=2.873787091e-16 puc=-2.202042248e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.042407714e+04 lvsat=-8.377842294e-03 wvsat=-7.743105575e-02 pvsat=3.045691929e-8 a0=1.051354951e+00 la0=1.721612128e-07 wa0=5.307471608e-07 pa0=-5.915185699e-13 ags=1.088237009e-01 lags=3.718389351e-07 wags=-6.002914877e-07 pags=8.644139931e-13 a1=0.0 a2=1.020591357e+00 la2=-2.181361750e-07 wa2=-1.267373402e-06 pa2=1.253267536e-12 b0=0.0 b1=0.0 keta=-1.316930213e-02 lketa=1.630631562e-09 wketa=8.978840231e-08 pketa=-9.917553844e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.388708941e-01 lpclm=-6.250535871e-08 wpclm=-3.075709197e-07 ppclm=4.461517458e-13 pdiblc1=1.308749221e+00 lpdiblc1=-8.955192397e-07 wpdiblc1=-4.729180260e-06 ppdiblc1=4.579666652e-12 pdiblc2=-1.595917611e-03 lpdiblc2=2.003369148e-09 wpdiblc2=4.420534383e-09 ppdiblc2=-4.371333835e-15 pdiblcb=1.172588168e-02 lpdiblcb=-3.631712262e-08 wpdiblcb=-1.853049166e-07 ppdiblcb=1.832424728e-13 drout=2.267188182e-01 ldrout=3.726861354e-08 wdrout=2.382882220e-06 pdrout=-1.699199387e-13 pscbe1=7.869784414e+08 lpscbe1=1.287662868e+01 wpscbe1=6.570186271e+01 ppscbe1=-6.497060098e-5 pscbe2=8.811227077e-09 lpscbe2=2.764390048e-16 wpscbe2=1.600634151e-15 ppscbe2=-9.896864416e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=7.058058197e-05 lalpha0=-3.450468022e-11 walpha0=-2.149614687e-10 palpha0=1.050882132e-16 alpha1=-3.989464227e-10 lalpha1=2.439199377e-16 walpha1=1.519602202e-15 palpha1=-7.428879284e-22 beta0=1.046580191e+02 lbeta0=-4.678903733e-05 wbeta0=-2.929793472e-04 pbeta0=1.437236978e-10 agidl=1.135120883e-08 lagidl=-5.748990419e-15 wagidl=-2.718830869e-14 pagidl=1.610640460e-20 bgidl=2.160768431e+09 lbgidl=-5.101142401e+02 wbgidl=-2.681233251e+03 pbgidl=1.427413095e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.924717974e-01 lkt1=6.351445455e-10 wkt1=1.169863187e-07 pkt1=-5.755947671e-14 kt2=-1.062481582e-01 lkt2=4.516400942e-08 wkt2=2.402369528e-07 pkt2=-1.676766103e-13 at=1.619462245e+05 lat=-4.275987261e-02 wat=2.091630816e-02 pat=-6.900685967e-8 ute=-6.913338111e+00 lute=3.258946807e-06 wute=2.111497117e-05 pute=-9.984413758e-12 ua1=-1.216904515e-08 lua1=7.442934724e-15 wua1=4.513708600e-14 pua1=-2.341278166e-20 ub1=7.951849306e-18 lub1=-5.015405048e-24 wub1=-2.741447983e-23 pub1=1.434568592e-29 uc1=8.020344020e-10 luc1=-5.642122732e-16 wuc1=-2.814004522e-15 puc1=1.795330719e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.009088881e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.262644252e-08 wvth0=-6.510265827e-08 pvth0=3.029418791e-14 k1=-1.602433399e-01 lk1=2.508268838e-07 wk1=1.912001661e-06 pk1=-6.127326464e-13 k2=2.443993654e-01 lk2=-8.619508927e-08 wk2=-7.071367771e-07 pk2=2.168561751e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.068204422e+00 ldsub=-3.334309579e-08 wdsub=9.969044353e-07 pdsub=-4.873566713e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.154691766e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.769023067e-08 wvoff=-2.698379294e-07 pvoff=7.111439303e-14 nfactor='3.890693957e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.407435114e-07 wnfactor=6.917066481e-06 pnfactor=-1.542716302e-12 eta0=-4.255318186e-01 leta0=2.186930855e-07 weta0=3.261040085e-07 peta0=-7.789646451e-14 etab=1.468804215e-03 letab=-5.001470127e-10 wetab=-5.631225722e-09 petab=1.345130888e-15 u0=6.817258769e-03 lu0=-7.344114957e-10 wu0=9.754171182e-09 pu0=-3.917054863e-16 ua=-1.740025874e-10 lua=-5.197311486e-16 wua=-2.372420517e-15 pua=1.267309373e-21 ub=-4.313896939e-19 lub=6.090516102e-25 wub=6.080935532e-24 pub=-1.912599479e-30 uc=4.643812610e-11 luc=-1.215541264e-17 wuc=-2.749743547e-16 puc=5.471331752e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.651255037e+04 lvsat=3.311785800e-03 wvsat=4.650700828e-02 pvsat=-3.013268208e-8 a0=2.079580100e+00 la0=-3.305072156e-07 wa0=-1.560859625e-06 pa0=4.310052396e-13 ags=2.600371964e-01 lags=2.979151935e-07 wags=8.649959848e-08 pags=5.286624347e-13 a1=0.0 a2=3.588172864e-01 la2=1.053853148e-07 wa2=2.534746804e-06 pa2=-6.054749690e-13 b0=0.0 b1=0.0 keta=1.248466783e-01 lketa=-6.584124079e-08 wketa=-4.641470125e-07 pketa=1.716268678e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=3.911359554e-01 lpclm=5.860482075e-08 wpclm=1.177023973e-06 ppclm=-2.796221592e-13 pdiblc1=-1.248307950e+00 lpdiblc1=3.545492998e-07 wpdiblc1=8.659583286e-06 ppdiblc1=-1.965698183e-12 pdiblc2=-4.006168681e-03 lpdiblc2=3.181668589e-09 wpdiblc2=-5.066483103e-09 ppdiblc2=2.665844032e-16 pdiblcb=-9.845176336e-02 lpdiblcb=1.754542271e-08 wpdiblcb=3.706098331e-07 ppdiblcb=-8.852757084e-14 drout=1.595081483e-01 ldrout=7.012589376e-08 wdrout=4.022714455e-06 pdrout=-9.715847233e-13 pscbe1=8.258287353e+08 lpscbe1=-6.116114504e+00 wpscbe1=-1.303220350e+02 ppscbe1=3.085960190e-5 pscbe2=2.922546860e-08 lpscbe2=-9.703471248e-15 wpscbe2=-6.059420221e-14 ppscbe2=2.941550321e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.927406842e+00 lbeta0=1.078709509e-08 wbeta0=2.723594253e-06 pbeta0=-8.365991510e-13 agidl=-2.215598056e-09 lagidl=8.834144642e-16 wagidl=1.400902077e-14 pagidl=-4.033733856e-21 bgidl=8.092245841e+08 lbgidl=1.506150006e+02 wbgidl=1.630286330e+03 pbgidl=-6.803594825e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.211002050e-01 lkt1=1.463071415e-08 wkt1=8.318063136e-08 pkt1=-4.103289036e-14 kt2=-2.863303573e-03 lkt2=-5.377744449e-09 wkt2=-1.295510512e-07 pkt2=1.310165126e-14 at=1.195361263e+05 lat=-2.202684788e-02 wat=-2.832856651e-01 pat=7.970835900e-8 ute=-4.180238036e-01 lute=8.358250165e-08 wute=1.154029435e-06 pute=-2.261081696e-13 ua1=5.600615966e-09 lua1=-1.244119505e-15 wua1=-9.425666971e-15 pua1=3.261311382e-21 ub1=-4.469482015e-18 lub1=1.057011195e-24 wub1=7.846933584e-24 pub1=-2.892561258e-30 uc1=-7.326917920e-10 luc1=1.860693213e-16 wuc1=2.154780101e-15 puc1=-6.337590194e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.204633568e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.768342149e-08 wvth0=3.986264031e-08 pvth0=5.221127037e-15 k1=1.123683124e+00 lk1=-5.586463061e-08 wk1=-3.467219483e-06 pk1=6.722019082e-13 k2=-1.730916407e-01 lk2=1.353098735e-08 wk2=1.094355253e-06 pk2=-2.134662261e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-8.515412636e-01 ldsub=4.252265561e-07 wdsub=4.552755307e-06 pdsub=-1.336742769e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.075863507e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.196673994e-08 wvoff=-4.151865636e-07 pvoff=1.058338213e-13 nfactor='2.054060570e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.979731058e-07 wnfactor=8.694250275e-07 pnfactor=-9.811618793e-14 eta0=0.49 etab=-0.000625 u0=-4.250043246e-03 lu0=1.909234937e-09 wu0=4.936687374e-08 pu0=-9.853991745e-15 ua=-5.413215412e-09 lua=7.317596187e-16 wua=1.619518404e-14 pua=-3.167934327e-21 ub=4.702947734e-18 lub=-6.173875712e-25 wub=-1.177555559e-23 pub=2.352780555e-30 uc=9.989659462e-11 luc=-2.492503702e-17 wuc=-4.460339370e-16 puc=9.557431995e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.139882183e+04 lvsat=4.533302136e-03 wvsat=-2.055026784e-01 pvsat=3.006487178e-8 a0=-3.102288004e-01 la0=2.403464363e-07 wa0=3.438720520e-06 pa0=-7.632444697e-13 ags=2.127753980e+00 lags=-1.482263147e-07 wags=7.847494198e-06 pags=-1.325206345e-12 a1=0.0 a2=1.697589778e+00 la2=-2.144072702e-07 wa2=-1.726210965e-06 pa2=4.123400132e-13 b0=0.0 b1=0.0 keta=-5.356557137e-01 lketa=9.193296559e-08 wketa=1.468935435e-06 pketa=-2.901285365e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=8.980595131e-01 lpclm=-6.248400946e-08 wpclm=-1.496372491e-06 ppclm=3.589720542e-13 pdiblc1=-8.579017139e-02 lpdiblc1=7.685867795e-08 wpdiblc1=7.914442929e-07 ppdiblc1=-8.623582152e-14 pdiblc2=1.321340355e-02 lpdiblc2=-9.315706302e-10 wpdiblc2=-2.951629803e-08 ppdiblc2=6.106911695e-15 pdiblcb=-2.732510397e-01 lpdiblcb=5.929972585e-08 wpdiblcb=2.222728831e-06 ppdiblcb=-5.309432359e-13 drout=1.503710032e+00 ldrout=-2.509636102e-07 wdrout=-5.052048418e-06 pdrout=1.196103884e-12 pscbe1=8.029075316e+08 lpscbe1=-6.409265698e-01 wpscbe1=-1.038654193e+01 ppscbe1=2.210610665e-6 pscbe2=-2.538909488e-08 lpscbe2=3.342309529e-15 wpscbe2=1.038486722e-13 ppscbe2=-9.864966207e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=7.949721164e+00 lbeta0=2.443268731e-07 wbeta0=6.501395521e-07 pbeta0=-3.413130265e-13 agidl=5.628622265e-09 lagidl=-9.903344440e-16 wagidl=-1.390809390e-14 pagidl=2.634827325e-21 bgidl=2.166143256e+09 lbgidl=-1.735121626e+02 wbgidl=-3.137448936e+03 pbgidl=4.585094407e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.241519049e+00 lkt1=1.867171635e-07 wkt1=2.246970569e-06 pkt1=-5.578973928e-13 kt2=5.724519438e-02 lkt2=-1.973586136e-08 wkt2=-3.345106921e-07 pkt2=6.206036067e-14 at=-4.108139137e+04 lat=1.633985856e-02 wat=5.085673676e-01 pat=-1.094415749e-7 ute=2.151349326e+00 lute=-5.301636579e-07 wute=-6.405249927e-06 pute=1.579576892e-12 ua1=2.175432288e-09 lua1=-4.259458801e-16 wua1=5.606891670e-15 pua1=-3.295159006e-22 ub1=-2.303763716e-18 lub1=5.396860653e-25 wub1=-4.543604880e-24 pub1=6.716666453e-32 uc1=1.183462596e-10 luc1=-1.721813812e-17 wuc1=-1.387329598e-15 puc1=2.123447243e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.042811398e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.216253229e-08 wvth0=-9.944270744e-08 pvth0=3.163941846e-14 k1=-8.773446680e-01 lk1=3.104425600e-07 wk1=3.635632938e-06 pk1=-5.803352740e-13 k2=5.282837761e-01 lk2=-1.154715083e-07 wk2=-1.099355141e-06 pk2=1.727892604e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.740083934e+00 ldsub=-1.314761622e-06 wdsub=-2.062615595e-05 pdsub=3.208692702e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.910698695e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.568696858e-08 wvoff=5.093841348e-07 pvoff=-5.536193319e-14 nfactor='7.149655223e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.292152873e-07 wnfactor=5.400140196e-06 pnfactor=-9.501174898e-13 eta0=1.893639354e+00 leta0=-2.608944467e-07 weta0=-2.169709277e-09 peta0=4.032838634e-16 etab=3.394336571e-01 letab=-6.320670259e-08 wetab=-1.038562351e-06 petab=1.930375841e-13 u0=2.339518169e-02 lu0=-3.036981957e-09 wu0=-4.674338824e-08 pu0=7.018029638e-15 ua=3.886184039e-09 lua=-9.230541356e-16 wua=-1.386346346e-14 pua=2.100153216e-21 ub=-2.266581811e-18 lub=6.158870009e-25 wub=1.035262472e-23 pub=-1.523331891e-30 uc=-2.384631360e-10 luc=3.545670372e-17 wuc=7.243663492e-16 puc=-1.123465953e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.415348850e+05 lvsat=-2.849222424e-02 wvsat=-8.251022740e-02 pvsat=1.023087012e-8 a0=3.048128637e+00 la0=-3.596759882e-07 wa0=-9.225689060e-06 pa0=1.513854164e-12 ags=1.25 a1=0.0 a2=-1.688871825e+00 la2=3.934501494e-07 wa2=5.608934900e-06 pa2=-9.095336286e-13 b0=0.0 b1=0.0 keta=7.688199399e-02 lketa=-1.266460429e-08 wketa=-1.444299522e-06 pketa=2.221474507e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=3.075543399e-02 lpclm=9.243158736e-08 wpclm=3.822085082e-06 ppclm=-5.934322421e-13 pdiblc1=1.572835776e+00 lpdiblc1=-2.236928288e-07 wpdiblc1=1.382822590e-06 ppdiblc1=-2.048365929e-13 pdiblc2=3.114521763e-02 lpdiblc2=-4.358337341e-09 wpdiblc2=3.613720176e-08 ppdiblc2=-5.481326679e-15 pdiblcb=-5.211727023e+00 lpdiblcb=9.831839101e-07 wpdiblcb=2.965908418e-05 ppdiblcb=-5.683988211e-12 drout=-5.086777361e+00 ldrout=9.487459873e-07 wdrout=1.258301368e-05 pdrout=-1.961314343e-12 pscbe1=7.944991595e+08 lpscbe1=8.574160031e-01 wpscbe1=1.675348074e+01 ppscbe1=-2.611365042e-6 pscbe2=-8.423568013e-08 lpscbe2=1.461659180e-14 wpscbe2=2.852497637e-13 ppscbe2=-4.457508489e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.566302834e+01 lbeta0=-1.164749353e-06 wbeta0=-6.104997183e-06 pbeta0=8.799045449e-13 agidl=-1.735479305e-09 lagidl=2.787349843e-16 wagidl=9.261134760e-15 pagidl=-1.406391369e-21 bgidl=8.467363718e+08 lbgidl=5.425867241e+01 wbgidl=4.667830778e+02 pbgidl=-1.652514064e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=1.108566154e+00 lkt1=-2.312965144e-07 wkt1=-3.052991049e-06 pkt1=3.710434147e-13 kt2=3.874109525e-01 lkt2=-8.309056328e-08 wkt2=-1.259690573e-06 pkt2=2.402711091e-13 at=-7.158538946e+04 lat=2.365455642e-02 wat=7.076571870e-02 pat=-3.908477318e-8 ute=-5.553492691e+00 lute=8.485642010e-07 wute=2.095135258e-05 pute=-3.346180148e-12 ua1=-1.307045851e-09 lua1=1.784627202e-16 wua1=1.346978432e-14 pua1=-1.824163845e-21 ub1=9.199194857e-19 lub1=-5.170191884e-27 wub1=-9.411370202e-24 pub1=9.786998163e-31 uc1=2.560730738e-11 luc1=-1.714084476e-18 wuc1=-1.590789406e-16 puc1=5.426338350e-24 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos lmin=2.0e-05 lmax=0.0001 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.143862851e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.103372644e-06 wvth0=8.837866606e-08 pvth0=-1.766589667e-12 k1=4.303698969e-01 lk1=1.109590230e-06 wk1=-1.863414147e-08 pk1=3.724754314e-13 k2=2.209900758e-02 lk2=-2.409044937e-07 wk2=3.082242674e-08 pk2=-6.161054813e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.121609426e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.498620184e-07 wvoff=-3.702486531e-08 pvoff=7.400852194e-13 nfactor='8.120382066e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.038328362e-06 wnfactor=-1.348751715e-06 pnfactor=2.696002270e-11 eta0=0.08 etab=-0.07 u0=3.513422016e-02 lu0=-4.416362437e-07 wu0=-4.229238861e-08 pu0=8.453770579e-13 ua=7.053534227e-10 lua=-2.629029356e-14 wua=-2.736587223e-15 pua=5.470128624e-20 ub=3.831042496e-18 lub=-4.327535737e-23 wub=-4.013641232e-24 pub=8.022815281e-29 uc=-6.496972548e-11 luc=-8.841609808e-16 wuc=-1.468731067e-17 puc=2.935827436e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.113870874e+05 lvsat=-3.019810289e+00 wvsat=-3.090414997e-01 pvsat=6.177390362e-6 a0=1.040300036e+00 la0=1.151561927e-05 wa0=1.317404103e-06 pa0=-2.633341935e-11 ags=3.874323218e-02 lags=8.789572236e-06 wags=9.715722784e-07 pags=-1.942063197e-11 a1=0.0 a2=1.561282690e+00 la2=-1.521718071e-05 wa2=-1.557296618e-06 pa2=3.112859965e-11 b0=0.0 b1=0.0 keta=8.574671297e-02 lketa=-2.338351742e-06 wketa=-2.875115450e-07 pketa=5.747030896e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.762746415e-01 lpclm=4.725784767e-06 wpclm=7.784550232e-07 ppclm=-1.556043626e-11 pdiblc1=0.39 pdiblc2=1.331171642e-02 lpdiblc2=-2.603495722e-07 wpdiblc2=-2.695201662e-08 ppdiblc2=5.387403565e-13 pdiblcb=7.855039219e-03 lpdiblcb=-1.876027773e-07 wpdiblcb=-2.312339226e-08 ppdiblcb=4.622104819e-13 drout=0.56 pscbe1=8.064388516e+08 lpscbe1=-3.234049569e+02 wpscbe1=-2.159460135e+02 ppscbe1=4.316516791e-3 pscbe2=9.285602072e-09 lpscbe2=1.497834542e-15 wpscbe2=7.781094574e-16 ppscbe2=-1.555352879e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-8.576215346e-10 lalpha0=1.914177236e-14 walpha0=2.916553213e-15 palpha0=-5.829860303e-20 alpha1=3.549704974e-10 lalpha1=-5.096572126e-15 walpha1=-7.765437562e-16 palpha1=1.552223219e-20 beta0=9.273771998e+00 lbeta0=-1.254056129e-04 wbeta0=-1.228462290e-05 pbeta0=2.455557302e-10 agidl=-9.457973221e-09 lagidl=1.940314624e-13 wagidl=3.123532565e-14 pagidl=-6.243588639e-19 bgidl=4.363286167e+08 lbgidl=1.126715400e+04 wbgidl=2.304639364e+03 pbgidl=-4.606713664e-2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.637968559e-01 lkt1=1.650452194e-07 wkt1=7.786872433e-08 pkt1=-1.556507808e-12 kt2=-0.037961 at=0.0 ute=-1.653904217e-01 lute=-3.284162913e-06 wute=-3.898887027e-07 pute=7.793434593e-12 ua1=2.139764998e-09 lua1=7.182700633e-15 ub1=-2.472812867e-19 lub1=-2.865441920e-23 wub1=-9.886991928e-25 pub1=1.976297963e-29 uc1=4.338507642e-11 luc1=7.645641303e-15 puc1=-3.308722450e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0886635+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.4858803 k2=0.010047076 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.64967492+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='8.0184089+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0130401126 ua=-6.0989319e-10 ub=1.66606982e-18 uc=-1.0920239e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160312.5 a0=1.6164016 ags=0.47846655 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-0.031235975 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.060146165 pdiblc1=0.39 pdiblc2=0.00028698955 pdiblcb=-0.0015303226 drout=0.56 pscbe1=790259600.0 pscbe2=9.3605355e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.0 agidl=2.4900183e-10 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.45554 kt2=-0.037961 at=0.0 ute=-0.32969 ua1=2.4991e-9 ub1=-1.6808e-18 uc1=4.2588e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.093883435e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.170138215e-8 k1=4.522972755e-01 lk1=2.682904169e-7 k2=2.243897693e-02 lk2=-9.899728555e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.724699858e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.821068169e-7 nfactor='8.375619887e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.853712138e-6 eta0=0.08 etab=-0.07 u0=1.610008706e-02 lu0=-2.444573819e-8 ua=-1.211989359e-10 lua=-3.904114865e-15 ub=1.642518584e-18 lub=1.881477614e-25 uc=-1.423307551e-10 luc=2.646582022e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.212579461e+05 lvsat=-4.868852462e-1 a0=1.673710294e+00 la0=-4.578317032e-7 ags=4.558541944e-01 lags=1.806471690e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-3.743565127e-02 lketa=4.952840774e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.109267259e-01 lpclm=4.562227086e-06 wpclm=1.110223025e-22 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=3.587787891e-04 lpdiblc2=-5.735148984e-10 pdiblcb=-4.459427061e-04 lpdiblcb=-8.662970003e-9 drout=0.56 pscbe1=7.805463027e+08 lpscbe1=7.759826970e+1 pscbe2=9.153007757e-09 lpscbe2=1.657912159e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-6.819567689e-01 lbeta0=2.941467397e-5 agidl=-4.042535850e-10 lagidl=5.218772587e-15 pagidl=1.654361225e-36 bgidl=8.022575536e+08 lbgidl=1.579738698e+3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.101376581e-01 lkt1=4.361735931e-7 kt2=-3.138933667e-02 lkt2=-5.250016399e-8 at=-1.789107917e+05 lat=1.429295056e+0 ute=1.617288118e-01 lute=-3.925881003e-6 ua1=5.328096354e-09 lua1=-2.260048410e-14 ub1=-4.224512371e-18 lub1=2.032138745e-23 uc1=7.901037197e-10 luc1=-2.909735948e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.091149793e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.079724093e-8 k1=5.977558582e-01 lk1=-3.119249599e-7 k2=-2.975396524e-02 lk2=1.091935757e-07 wk2=3.469446952e-24 pk2=-6.938893904e-30 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.915414784e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.581805218e-7 nfactor='8.421149226e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.035322754e-6 eta0=0.08 etab=-0.07 u0=8.149894523e-03 lu0=7.266546324e-9 ua=-1.665485757e-09 lua=2.255844507e-15 ub=2.098150966e-18 lub=-1.629310578e-24 uc=-6.694967090e-11 luc=-3.602714318e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.447013512e+05 lvsat=-1.815109412e-1 a0=1.964587897e+00 la0=-1.618104650e-6 ags=6.476342087e-01 lags=-5.843383766e-07 wags=-8.881784197e-22 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-4.118284482e-02 lketa=6.447547569e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.336218480e-01 lpclm=-1.199889384e-6 pdiblc1=0.39 pdiblc2=0.000215 pdiblcb=1.963998626e-02 lpdiblcb=-8.878312947e-08 wpdiblcb=-6.938893904e-24 ppdiblcb=1.387778781e-29 drout=0.56 pscbe1=800000000.0 pscbe2=1.671893803e-08 lpscbe2=-2.852160011e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.565947440e+00 lbeta0=4.492596311e-6 agidl=5.125510518e-10 lagidl=1.561758076e-15 bgidl=1.143013757e+09 lbgidl=2.205064997e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.434839429e-01 lkt1=-2.285864121e-7 kt2=-4.017360155e-02 lkt2=-1.746087337e-8 at=2.745973838e+05 lat=-3.796900997e-1 ute=-1.640382899e+00 lute=3.262508336e-6 ua1=-3.274541222e-09 lua1=1.171431885e-14 wua1=-8.271806126e-31 pua1=-1.654361225e-36 ub1=3.170152177e-18 lub1=-9.174968124e-24 uc1=9.216446460e-11 luc1=-1.257469911e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.090845143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.019133174e-8 k1=4.322967437e-01 lk1=1.715170913e-8 k2=2.844424485e-02 lk2=-6.555098444e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.916658762e-01 ldsub=3.347946888e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.722230050e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.087158959e-8 nfactor='8.494631950e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.181470339e-6 eta0=-5.744849986e-02 leta0=2.733671979e-07 peta0=1.110223025e-28 etab=6.842919891e-01 letab=-1.500188708e-06 wetab=-3.330669074e-22 petab=-1.110223025e-28 u0=1.359424468e-02 lu0=-3.561558378e-9 ua=-1.917591780e-10 lua=-6.752060745e-16 ub=1.151418582e-18 lub=2.536170597e-25 uc=-1.214437714e-10 luc=7.235453841e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.038194939e+04 lvsat=2.596678738e-2 a0=1.099283968e+00 la0=1.028723755e-7 ags=1.353546988e-01 lags=4.345189724e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-2.629453859e-03 lketa=-1.220220699e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.108255342e-02 lpclm=5.752552428e-7 pdiblc1=4.088045794e-01 lpdiblc1=-3.739986375e-8 pdiblc2=2.392950000e-06 lpdiblc2=4.228477835e-10 pdiblcb=-0.025 drout=1.344068365e-01 ldrout=8.464494752e-7 pscbe1=800000000.0 pscbe2=-4.454152232e-09 lpscbe2=1.358892391e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.794355910e+00 lbeta0=2.049451557e-6 agidl=6.445524780e-10 lagidl=1.299224399e-15 bgidl=1.269088568e+09 lbgidl=-3.023991007e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.444605805e-01 lkt1=-2.775700689e-8 kt2=-6.040588351e-02 lkt2=2.277850526e-8 at=6.493100483e+04 lat=3.730907145e-2 ute=0.0 ua1=2.824339679e-09 lua1=-4.155624112e-16 ub1=-1.527062104e-18 lub1=1.671804431e-25 uc1=1.528486051e-10 luc1=-2.464398577e-16 wuc1=-5.169878828e-32 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.084139568e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.356038974e-8 k1=3.328536151e-01 lk1=1.154880357e-7 k2=6.118412774e-02 lk2=-3.893058644e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=4.664626476e-01 ldsub=2.608304055e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.014237749e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.974735493e-8 nfactor='5.907109181e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.227466980e-7 eta0=3.582529886e-01 leta0=-1.377075330e-7 etab=-1.646537114e+00 letab=8.046982669e-7 u0=1.169191212e-02 lu0=-1.680398776e-9 ua=-5.906662208e-10 lua=-2.807388671e-16 ub=1.291920204e-18 lub=1.146792206e-25 uc=-6.422249855e-11 luc=1.577013837e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.500035228e+04 lvsat=1.622387311e-3 a0=1.225620556e+00 la0=-2.205808617e-8 ags=-8.827609932e-02 lags=6.556607597e-07 pags=4.440892099e-28 a1=0.0 a2=6.044617774e-01 la2=1.933618822e-7 b0=0.0 b1=0.0 keta=1.631183582e-02 lketa=-3.093268012e-08 pketa=-1.387778781e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.378830106e-01 lpclm=8.398417474e-8 pdiblc1=-2.440305587e-01 lpdiblc1=6.081692192e-7 pdiblc2=-1.444786656e-04 lpdiblc2=5.680847180e-10 pdiblcb=-4.911716338e-02 lpdiblcb=2.384873935e-8 drout=1.009114736e+00 ldrout=-1.852292549e-8 pscbe1=8.085510012e+08 lpscbe1=-8.455828520e+0 pscbe2=9.336779542e-09 lpscbe2=-4.851479500e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.461134792e+00 lbeta0=4.012239235e-7 agidl=2.424195336e-09 lagidl=-4.606110339e-16 bgidl=1.280411890e+09 lbgidl=-4.143720287e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.540604914e-01 lkt1=-1.826394297e-8 kt2=-2.736871980e-02 lkt2=-9.890954821e-9 at=1.688138884e+05 lat=-6.541759562e-2 ute=1.955480000e-02 lute=-1.933715508e-8 ua1=2.651272672e-09 lua1=-2.444216402e-16 wua1=-3.308722450e-30 ub1=-1.049425256e-18 lub1=-3.051403071e-25 uc1=-1.219162794e-10 luc1=2.526689368e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.030464698e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.679644165e-9 k1=4.675435820e-01 lk1=4.964215164e-8 k2=1.221796632e-02 lk2=-1.499249910e-08 pk2=6.938893904e-30 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.395528179e+00 ldsub=-1.933618609e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.040678042e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.103994151e-8 nfactor='6.161844639e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.472792213e-07 wnfactor=-7.105427358e-21 eta0=-3.184587778e-01 leta0=1.931165483e-07 peta0=5.551115123e-29 etab=-3.801533128e-04 letab=-5.848652817e-11 u0=1.001994485e-02 lu0=-8.630241358e-10 ua=-9.529635079e-10 lua=-1.036225924e-16 ub=1.565225622e-18 lub=-1.893159938e-26 uc=-4.384699617e-11 luc=5.809166520e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.178266868e+04 lvsat=-6.581983708e-3 a0=1.567087208e+00 la0=-1.889908884e-7 ags=2.884384880e-01 lags=4.714962994e-7 a1=0.0 a2=1.191076445e+00 la2=-9.341643046e-8 b0=0.0 b1=0.0 keta=-2.755142380e-02 lketa=-9.489248387e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=7.776001892e-01 lpclm=-3.320636238e-8 pdiblc1=1.594980969e+00 lpdiblc1=-2.908683466e-7 pdiblc2=-5.669698530e-03 lpdiblc2=3.269198953e-9 pdiblcb=2.323432675e-02 lpdiblcb=-1.152173363e-08 wpdiblcb=-9.540979118e-24 ppdiblcb=-6.396792818e-30 drout=1.480326837e+00 ldrout=-2.488843850e-7 pscbe1=7.830387781e+08 lpscbe1=4.016331970e+0 pscbe2=9.329958843e-09 lpscbe2=-4.518035983e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=9.821672202e+00 lbeta0=-2.639019999e-7 agidl=2.384125997e-09 lagidl=-4.410223361e-16 bgidl=1.344513051e+09 lbgidl=-7.277433743e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.937886636e-01 lkt1=1.157968567e-9 kt2=-4.540011584e-02 lkt2=-1.075946241e-9 at=2.652206705e+04 lat=4.144607083e-3 ute=-3.910960000e-02 lute=9.342110152e-9 ua1=2.505791010e-09 lua1=-1.733000203e-16 ub1=-1.893018625e-18 lub1=1.072671831e-25 uc1=-2.519095944e-11 luc1=-2.201921350e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.073748297e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.596912098e-08 wvth0=-6.569670674e-14 pvth0=1.569297314e-20 k1=-1.474413380e-02 lk1=1.648462183e-07 wk1=-3.816552709e-13 pk1=9.116599431e-20 k2=1.862291287e-01 lk2=-5.655854547e-08 wk2=1.250127735e-14 pk2=-2.986180192e-21 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=6.433110956e-01 ldsub=-1.367976616e-08 wdsub=7.455866324e-14 pdsub=-1.780982783e-20 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.439087585e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.278275029e-08 wvoff=-3.922896319e-14 pvoff=9.370622722e-21 nfactor='2.339527582e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.657576542e-07 wnfactor=4.173395070e-13 pnfactor=-9.968988834e-20 eta0=0.49 etab=-0.000625 u0=1.195908546e-02 lu0=-1.326226653e-09 wu0=-5.246282853e-15 pu0=1.253179588e-21 ua=-9.568609602e-11 lua=-3.084004478e-16 wua=-2.315927408e-22 pua=5.532055806e-29 ub=8.365600827e-19 lub=1.551247380e-25 wub=-2.955879191e-31 pub=7.060708546e-38 uc=-4.655425743e-11 luc=6.455850017e-18 wuc=-7.089599594e-26 puc=1.693493330e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.075953780e+03 lvsat=1.440480544e-02 wvsat=-1.737638842e-08 pvsat=4.150697903e-15 a0=8.188412249e-01 la0=-1.025737040e-08 wa0=1.110700154e-14 pa0=-2.653129272e-21 ags=4.704401308e+00 lags=-5.833447395e-07 wags=4.100134916e-13 pags=-9.793992106e-20 a1=0.0 a2=1.130805108e+00 la2=-7.901941609e-08 wa2=8.951765587e-13 pa2=-2.138308242e-19 b0=0.0 b1=0.0 keta=-5.334522481e-02 lketa=-3.327883141e-09 wketa=-5.907980771e-16 pketa=1.411240014e-22 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.067403384e-01 lpclm=5.538093019e-08 wpclm=-3.899264911e-15 ppclm=9.314176097e-22 pdiblc1=1.740727862e-01 lpdiblc1=4.854399118e-08 wpdiblc1=-4.785460561e-14 ppdiblc1=1.143102946e-20 pdiblc2=3.522017863e-03 lpdiblc2=1.073573658e-09 wpdiblc2=-5.742553377e-16 ppdiblc2=1.371723707e-22 pdiblcb=4.565600017e-01 lpdiblcb=-1.150302376e-07 wpdiblcb=2.677494785e-13 ppdiblcb=-6.395731800e-20 drout=-1.550803608e-01 ldrout=1.417653322e-07 wdrout=9.618185182e-14 pdrout=-2.297495882e-20 pscbe1=7.994972153e+08 lpscbe1=8.490506716e-02 wpscbe1=-7.798528671e-06 ppscbe1=1.862834930e-12 pscbe2=8.708594014e-09 lpscbe2=1.032450570e-16 wpscbe2=7.999399536e-22 ppscbe2=-1.910816596e-28 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.163187944e+00 lbeta0=1.322601349e-07 wbeta0=4.312823023e-13 pbeta0=-1.030204047e-19 agidl=1.062036611e-09 lagidl=-1.252148444e-16 wagidl=-1.666049370e-22 pagidl=3.979692113e-29 bgidl=1.135992664e+09 lbgidl=-2.296507275e+01 wbgidl=3.698393135e-04 pbgidl=-8.834351635e-11 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.037483494e-01 lkt1=3.537038708e-09 wkt1=-1.061072474e-13 pkt1=2.534583832e-20 kt2=-5.258809566e-02 lkt2=6.410464987e-10 wkt2=-7.603565111e-15 pkt2=1.816263584e-21 at=1.259016779e+05 lat=-1.959420056e-02 wat=5.825264635e-08 pat=-1.391480965e-14 ute=4.824857555e-02 lute=-1.152513724e-08 wute=-1.254854221e-14 pute=2.997470272e-21 ua1=4.016400244e-09 lua1=-5.341392479e-16 wua1=-8.401142233e-22 pua1=2.006780839e-28 ub1=-3.795611892e-18 lub1=5.617396367e-25 wub1=7.444050248e-31 pub1=-1.778160289e-37 uc1=-3.371697339e-10 luc1=5.250315636e-17 wuc1=-6.676013217e-23 puc1=1.594699272e-29 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.075462027e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.177411773e-08 wvth0=-1.234542140e-12 pvth0=2.345260706e-19 k1=3.163794938e-01 lk1=1.198951989e-07 wk1=3.685256118e-13 pk1=-3.909252211e-20 k2=1.673213808e-01 lk2=-5.873786326e-08 wk2=-1.282034932e-13 pk2=2.286599943e-20 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.967688838e+00 ldsub=-2.612189876e-07 wdsub=-4.483775840e-13 pdsub=7.759543186e-20 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.238186134e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.750942367e-08 wvoff=2.986523207e-14 pvoff=-2.528583121e-21 nfactor='8.922740736e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.041177492e-06 wnfactor=-8.050367853e-12 pnfactor=1.464167187e-18 eta0=1.892926871e+00 leta0=-2.607620175e-07 weta0=2.447968441e-13 peta0=-4.550038968e-20 etab=-1.568066564e-03 letab=1.752877822e-10 wetab=8.391869422e-16 petab=-1.559796775e-22 u0=8.047446303e-03 lu0=-7.326803986e-10 wu0=1.230471539e-14 pu0=-1.882867928e-21 ua=-6.657480479e-10 lua=-2.334894449e-16 wua=1.045366863e-21 pua=-1.764588485e-28 ub=1.132600365e-18 lub=1.157160070e-25 wub=7.047681971e-31 pub=-1.082211513e-37 uc=-6.245784946e-13 luc=-1.431194449e-18 wuc=6.015200804e-24 puc=-1.112583075e-30 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.144435132e+05 lvsat=-2.513302832e-02 wvsat=-1.495893276e-07 pvsat=2.914296417e-14 a0=1.896421654e-02 la0=1.373831684e-07 wa0=7.414769492e-13 pa0=-1.386740793e-19 ags=1.250000346e+00 lags=-5.389125057e-14 wags=-1.053008134e-12 pags=1.641323779e-19 a1=0.0 a2=1.527674086e-01 la2=9.481363330e-08 wa2=-2.065570250e-12 pa2=3.149570160e-19 b0=0.0 b1=0.0 keta=-3.973396729e-01 lketa=6.027534974e-08 wketa=4.199554233e-13 pketa=-7.801159535e-20 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.285699180e+00 lpclm=-1.024159983e-07 wpclm=8.004728080e-13 ppclm=-1.484834549e-19 pdiblc1=2.026872356e+00 lpdiblc1=-2.909489823e-07 wpdiblc1=-1.206082928e-12 ppdiblc1=2.278616802e-19 pdiblc2=4.301049316e-02 lpdiblc2=-6.158073494e-09 wpdiblc2=5.757148719e-14 ppdiblc2=-1.065656776e-20 pdiblcb=4.526545287e+00 lpdiblcb=-8.830983993e-07 wpdiblcb=-1.221049108e-11 ppdiblcb=2.248934727e-18 drout=-9.552692295e-01 ldrout=3.047678332e-07 wdrout=1.623279807e-12 pdrout=-3.091295264e-19 pscbe1=7.999999934e+08 lpscbe1=1.025021076e-06 wpscbe1=2.002840424e-05 ppscbe1=-3.121827126e-12 pscbe2=9.423272207e-09 lpscbe2=-1.919858632e-17 wpscbe2=-1.991224164e-21 ppscbe2=3.084759924e-28 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.365851252e+01 lbeta0=-8.758413281e-07 wbeta0=3.080038482e-13 pbeta0=-9.047761296e-20 agidl=1.305323381e-09 lagidl=-1.830398288e-16 wagidl=-7.961726653e-22 pagidl=1.608209977e-28 bgidl=1.000000312e+09 lbgidl=-4.861084700e-05 wbgidl=-9.498316803e-04 pbgidl=1.480502644e-10 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.061462833e-01 lkt1=-1.094680060e-07 wkt1=9.623834067e-13 pkt1=-1.707029753e-19 kt2=-2.619607966e-02 lkt2=-4.199903906e-09 wkt2=1.035279331e-13 pkt2=-1.865690624e-20 at=-4.835015559e+04 lat=1.082145614e-02 wat=-2.075133112e-08 pat=-6.311324396e-16 ute=1.325677818e+00 lute=-2.501211363e-07 wute=-4.604924002e-13 pute=8.655854808e-20 ua1=3.115624181e-09 lua1=-4.204833471e-16 wua1=3.175666108e-21 pua1=-5.255329125e-28 ub1=-2.170210357e-18 lub1=3.161761073e-25 wub1=-2.771513092e-30 pub1=4.577870828e-37 uc1=-2.662475279e-11 luc1=6.760904313e-20 wuc1=1.709455309e-22 puc1=-2.662998859e-29 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos lmin=2.0e-05 lmax=0.0001 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.100659040e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.397772846e-7 k1=4.212606180e-01 lk1=1.291674424e-6 k2=3.716651602e-02 lk2=-5.420869610e-7 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.302605061e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.880721963e-7 nfactor='7.461046316e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.114104823e-5 eta0=0.08 etab=-0.07 u0=1.445963384e-02 lu0=-2.837462552e-8 ua=-6.324241445e-10 lua=4.503683210e-16 ub=1.868978521e-18 lub=-4.055915651e-24 wub=-3.081487911e-39 uc=-7.214960068e-11 luc=-7.406433888e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160312.5 a0=1.684311541e+00 la0=-1.357442978e-6 ags=5.136952411e-01 lags=-7.041817269e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-5.480298045e-02 lketa=4.710778082e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.042722157e-01 lpclm=-2.880916892e-6 pdiblc1=0.39 pdiblc2=1.362535913e-04 lpdiblc2=3.013041483e-9 pdiblcb=-3.448804924e-03 lpdiblcb=3.834829377e-8 drout=0.56 pscbe1=7.008738872e+08 lpscbe1=1.786719392e+3 pscbe2=9.665980000e-09 lpscbe2=-6.105490408e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=5.681322036e-10 lalpha0=-9.357433760e-15 alpha1=-2.464203913e-11 lalpha1=2.491453517e-15 palpha1=-2.197198502e-37 beta0=3.268447993e+00 lbeta0=-5.365972042e-6 agidl=5.811380381e-09 lagidl=-1.111856617e-13 bgidl=1.562948962e+09 lbgidl=-1.125271361e+4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.257308181e-01 lkt1=-5.958518612e-7 kt2=-0.037961 at=0.0 ute=-3.559870728e-01 lute=5.256487698e-7 ua1=2.139764998e-09 lua1=7.182700633e-15 ub1=-7.306057684e-19 lub1=-1.899330897e-23 uc1=4.338507642e-11 luc1=7.645641303e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0886635+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.4858803 k2=0.010047076 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.64967492+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='8.0184089+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0130401126 ua=-6.0989319e-10 ub=1.66606982e-18 uc=-1.0920239e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160312.5 a0=1.6164016 ags=0.47846655 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-0.031235975 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.060146165 pdiblc1=0.39 pdiblc2=0.00028698955 pdiblcb=-0.0015303226 drout=0.56 pscbe1=790259600.0 pscbe2=9.3605355e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.0 agidl=2.4900183e-10 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.45554 kt2=-0.037961 at=0.0 ute=-0.32969 ua1=2.4991e-9 ub1=-1.6808e-18 uc1=4.2588e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.093883435e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.170138215e-8 k1=4.522972755e-01 lk1=2.682904169e-7 k2=2.243897693e-02 lk2=-9.899728555e-08 pk2=1.110223025e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.724699858e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.821068169e-7 nfactor='8.375619887e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.853712138e-6 eta0=0.08 etab=-0.07 u0=1.610008706e-02 lu0=-2.444573819e-8 ua=-1.211989359e-10 lua=-3.904114865e-15 ub=1.642518584e-18 lub=1.881477614e-25 uc=-1.423307551e-10 luc=2.646582022e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.212579461e+05 lvsat=-4.868852462e-1 a0=1.673710294e+00 la0=-4.578317032e-7 ags=4.558541944e-01 lags=1.806471690e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-3.743565127e-02 lketa=4.952840774e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.109267259e-01 lpclm=4.562227086e-06 wpclm=-4.440892099e-22 pdiblc1=0.39 pdiblc2=3.587787891e-04 lpdiblc2=-5.735148984e-10 pdiblcb=-4.459427061e-04 lpdiblcb=-8.662970003e-9 drout=0.56 pscbe1=7.805463027e+08 lpscbe1=7.759826970e+1 pscbe2=9.153007757e-09 lpscbe2=1.657912159e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-6.819567689e-01 lbeta0=2.941467397e-5 agidl=-4.042535850e-10 lagidl=5.218772587e-15 bgidl=8.022575536e+08 lbgidl=1.579738698e+3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.101376581e-01 lkt1=4.361735931e-7 kt2=-3.138933667e-02 lkt2=-5.250016399e-8 at=-1.789107917e+05 lat=1.429295056e+0 ute=1.617288118e-01 lute=-3.925881003e-6 ua1=5.328096354e-09 lua1=-2.260048410e-14 pua1=-2.646977960e-35 ub1=-4.224512371e-18 lub1=2.032138745e-23 pub1=2.465190329e-44 uc1=7.901037197e-10 luc1=-2.909735948e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.091149793e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.079724093e-8 k1=5.977558582e-01 lk1=-3.119249599e-7 k2=-2.975396524e-02 lk2=1.091935757e-07 wk2=2.081668171e-23 pk2=-1.387778781e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.915414784e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.581805218e-7 nfactor='8.421149226e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.035322754e-6 eta0=0.08 etab=-0.07 u0=8.149894523e-03 lu0=7.266546324e-9 ua=-1.665485757e-09 lua=2.255844507e-15 ub=2.098150966e-18 lub=-1.629310578e-24 uc=-6.694967090e-11 luc=-3.602714318e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.447013512e+05 lvsat=-1.815109412e-1 a0=1.964587897e+00 la0=-1.618104650e-6 ags=6.476342087e-01 lags=-5.843383766e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-4.118284482e-02 lketa=6.447547569e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.336218480e-01 lpclm=-1.199889384e-06 wpclm=1.776356839e-21 pdiblc1=0.39 pdiblc2=0.000215 pdiblcb=1.963998626e-02 lpdiblcb=-8.878312947e-08 ppdiblcb=-4.163336342e-29 drout=0.56 pscbe1=800000000.0 pscbe2=1.671893803e-08 lpscbe2=-2.852160011e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.565947440e+00 lbeta0=4.492596311e-6 agidl=5.125510518e-10 lagidl=1.561758076e-15 bgidl=1.143013757e+09 lbgidl=2.205064997e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.434839429e-01 lkt1=-2.285864121e-7 kt2=-4.017360155e-02 lkt2=-1.746087337e-8 at=2.745973838e+05 lat=-3.796900997e-1 ute=-1.640382899e+00 lute=3.262508336e-6 ua1=-3.274541222e-09 lua1=1.171431885e-14 wua1=8.271806126e-31 pua1=8.271806126e-36 ub1=3.170152177e-18 lub1=-9.174968124e-24 wub1=3.081487911e-39 pub1=6.162975822e-45 uc1=9.216446460e-11 luc1=-1.257469911e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.090845143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.019133174e-8 k1=4.322967437e-01 lk1=1.715170913e-8 k2=2.844424485e-02 lk2=-6.555098444e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.916658762e-01 ldsub=3.347946888e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.722230050e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.087158959e-8 nfactor='8.494631950e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.181470339e-6 eta0=-5.744849986e-02 leta0=2.733671979e-7 etab=6.842919891e-01 letab=-1.500188708e-06 wetab=2.220446049e-22 petab=-1.554312234e-27 u0=1.359424468e-02 lu0=-3.561558378e-9 ua=-1.917591780e-10 lua=-6.752060745e-16 ub=1.151418582e-18 lub=2.536170597e-25 uc=-1.214437714e-10 luc=7.235453841e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.038194939e+04 lvsat=2.596678738e-2 a0=1.099283968e+00 la0=1.028723755e-7 ags=1.353546988e-01 lags=4.345189724e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-2.629453859e-03 lketa=-1.220220699e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.108255342e-02 lpclm=5.752552428e-7 pdiblc1=4.088045794e-01 lpdiblc1=-3.739986375e-8 pdiblc2=2.392950000e-06 lpdiblc2=4.228477835e-10 pdiblcb=-0.025 drout=1.344068365e-01 ldrout=8.464494752e-7 pscbe1=800000000.0 pscbe2=-4.454152232e-09 lpscbe2=1.358892391e-14 ppscbe2=1.323488980e-35 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.794355910e+00 lbeta0=2.049451557e-6 agidl=6.445524780e-10 lagidl=1.299224399e-15 bgidl=1.269088568e+09 lbgidl=-3.023991007e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.444605805e-01 lkt1=-2.775700689e-8 kt2=-6.040588351e-02 lkt2=2.277850526e-8 at=6.493100483e+04 lat=3.730907145e-2 ute=0.0 ua1=2.824339679e-09 lua1=-4.155624112e-16 ub1=-1.527062104e-18 lub1=1.671804431e-25 uc1=1.528486051e-10 luc1=-2.464398577e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.084139568e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.356038974e-8 k1=3.328536151e-01 lk1=1.154880357e-7 k2=6.118412774e-02 lk2=-3.893058644e-08 pk2=2.775557562e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=4.664626476e-01 ldsub=2.608304055e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.014237749e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.974735493e-8 nfactor='5.907109181e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.227466980e-7 eta0=3.582529886e-01 leta0=-1.377075330e-7 etab=-1.646537114e+00 letab=8.046982669e-7 u0=1.169191212e-02 lu0=-1.680398776e-9 ua=-5.906662208e-10 lua=-2.807388671e-16 ub=1.291920204e-18 lub=1.146792206e-25 uc=-6.422249855e-11 luc=1.577013837e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.500035228e+04 lvsat=1.622387311e-3 a0=1.225620556e+00 la0=-2.205808617e-8 ags=-8.827609932e-02 lags=6.556607597e-7 a1=0.0 a2=6.044617774e-01 la2=1.933618822e-7 b0=0.0 b1=0.0 keta=1.631183582e-02 lketa=-3.093268012e-08 pketa=-2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.378830106e-01 lpclm=8.398417474e-8 pdiblc1=-2.440305587e-01 lpdiblc1=6.081692192e-7 pdiblc2=-1.444786656e-04 lpdiblc2=5.680847180e-10 pdiblcb=-4.911716338e-02 lpdiblcb=2.384873935e-8 drout=1.009114736e+00 ldrout=-1.852292549e-8 pscbe1=8.085510012e+08 lpscbe1=-8.455828520e+0 pscbe2=9.336779542e-09 lpscbe2=-4.851479500e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.461134792e+00 lbeta0=4.012239235e-7 agidl=2.424195336e-09 lagidl=-4.606110339e-16 bgidl=1.280411890e+09 lbgidl=-4.143720287e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.540604914e-01 lkt1=-1.826394297e-8 kt2=-2.736871980e-02 lkt2=-9.890954821e-9 at=1.688138884e+05 lat=-6.541759562e-2 ute=1.955480000e-02 lute=-1.933715508e-8 ua1=2.651272672e-09 lua1=-2.444216402e-16 ub1=-1.049425256e-18 lub1=-3.051403071e-25 uc1=-1.219162794e-10 luc1=2.526689368e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.530901967e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.419691234e-07 wvth0=1.023705487e-06 pvth0=-5.004589013e-13 k1=1.941485345e+00 lk1=-6.709237583e-07 wk1=-3.015127698e-06 pk1=1.474005478e-12 k2=-4.934896120e-01 lk2=2.322327647e-07 wk2=1.034486548e-06 pk2=-5.057294386e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.273213053e+00 ldsub=-1.335656650e-07 wdsub=2.502105136e-07 pdsub=-1.223204138e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.897732128e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.835255362e-09 wvoff=-2.338035306e-07 pvoff=1.142995320e-13 nfactor='7.643935000e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.471828736e-06 wnfactor=-3.031796649e-06 pnfactor=1.482154428e-12 eta0=-3.184587778e-01 leta0=1.931165483e-07 weta0=2.220446049e-22 peta0=2.220446049e-28 etab=-3.801533128e-04 letab=-5.848652817e-11 u0=-1.838255122e-03 lu0=4.934094083e-09 wu0=2.425739474e-08 pu0=-1.185871257e-14 ua=-3.710467694e-09 lua=1.244438479e-15 wua=5.640811229e-15 pua=-2.757623385e-21 ub=2.952244514e-18 lub=-6.970035250e-25 wub=-2.837316359e-24 pub=1.387078849e-30 uc=1.387676902e-11 luc=-2.241025057e-17 wuc=-1.180810040e-16 puc=5.772626043e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.105805374e+05 lvsat=-6.954739778e-02 wvsat=-2.634717538e-01 pvsat=1.288034363e-7 a0=1.475372854e+00 la0=-1.441544921e-07 wa0=1.876129005e-07 pa0=-9.171831865e-14 ags=-4.927428888e+00 lags=3.021377384e-06 wags=1.066969305e-05 pags=-5.216092843e-12 a1=0.0 a2=4.845383075e-01 la2=2.519888689e-07 wa2=1.445309958e-06 pa2=-7.065686794e-13 b0=0.0 b1=0.0 keta=-5.730706253e-02 lketa=5.057390717e-09 wketa=6.086878920e-08 pketa=-2.975692498e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.272778334e+00 lpclm=-2.752841019e-07 wpclm=-1.012947306e-06 ppclm=4.951995497e-13 pdiblc1=2.029027959e+00 lpdiblc1=-5.030608985e-07 wpdiblc1=-8.878960716e-07 ppdiblc1=4.340657525e-13 pdiblc2=3.929458420e-03 lpdiblc2=-1.423540905e-09 wpdiblc2=-1.963624664e-08 ppdiblc2=9.599571893e-15 pdiblcb=-1.005287123e+00 lpdiblcb=4.912915477e-07 wpdiblcb=2.103966106e-06 ppdiblcb=-1.028565910e-12 drout=2.747894712e+00 ldrout=-8.685602921e-07 wdrout=-2.592964732e-06 pdrout=1.267622668e-12 pscbe1=7.837979489e+08 lpscbe1=3.645196149e+00 wpscbe1=-1.552976458e+00 ppscbe1=7.592036010e-7 pscbe2=1.025310421e-08 lpscbe2=-4.964784350e-16 wpscbe2=-1.888406470e-15 ppscbe2=9.231852710e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.100425080e+01 lbeta0=-8.420291984e-07 wbeta0=-2.419108794e-06 pbeta0=1.182629716e-12 agidl=1.264541260e-09 lagidl=1.063090545e-16 wagidl=2.290247169e-15 pagidl=-1.119633134e-21 bgidl=1.139174799e+09 lbgidl=2.760937388e+01 wbgidl=4.200444459e+02 pbgidl=-2.053471283e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.621627884e-01 lkt1=-1.430297303e-08 wkt1=-6.469458603e-08 pkt1=3.162724227e-14 kt2=-3.966831155e-02 lkt2=-3.878053400e-09 wkt2=-1.172510494e-08 pkt2=5.732052052e-15 at=-1.486758419e+05 lat=8.979360882e-02 wat=3.583886969e-01 pat=-1.752054822e-7 ute=-1.421594275e-01 lute=5.972007931e-08 wute=2.108009942e-07 pute=-1.030542820e-13 ua1=-2.270113440e-09 lua1=2.161496388e-15 wua1=9.769695213e-15 pua1=-4.776110899e-21 ub1=3.129669595e-18 lub1=-2.348174407e-24 wub1=-1.027452152e-23 pub1=5.022905337e-30 uc1=4.442561789e-10 luc1=-2.515178360e-16 wuc1=-9.603113940e-16 puc1=4.694674312e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='9.799010983e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.577864047e-07 wvth0=-3.656091024e-06 pvth0=6.174040912e-13 k1=-5.278822047e+00 lk1=1.053791069e-06 wk1=1.076831321e-05 pk1=-1.818445051e-12 k2=1.992327629e+00 lk2=-3.615543996e-07 wk2=-3.694594814e-06 pk2=6.239062262e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.080150869e+00 ldsub=-8.744890130e-08 wdsub=-8.936089771e-07 pdsub=1.509037480e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.521037468e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=8.171463930e-08 wvoff=8.350126091e-07 pvoff=-1.410085793e-13 nfactor='-2.953652076e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.059616889e-06 wnfactor=1.082784517e-05 pnfactor=-1.828498215e-12 eta0=0.49 etab=-0.000625 u0=5.430979707e-02 lu0=-8.477991144e-09 wu0=-8.663355264e-08 pu0=1.462980803e-14 ua=9.752543028e-09 lua=-1.971470892e-15 wua=-2.014575439e-14 pua=3.402013544e-21 ub=-4.117078961e-18 lub=9.916457734e-25 wub=1.013327271e-23 pub=-1.711205763e-30 uc=-2.527105617e-10 luc=4.126946513e-17 wuc=4.217178714e-16 puc=-7.121549695e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.660683505e+05 lvsat=9.208372207e-02 wvsat=9.409705492e-01 pvsat=-1.589016967e-7 a0=1.146392495e+00 la0=-6.557095375e-08 wa0=-6.700460731e-07 pa0=1.131506804e-13 ags=2.333249928e+01 lags=-3.729071658e-06 wags=-3.810604662e-05 pags=6.434968093e-12 a1=0.0 a2=3.654156037e+00 la2=-5.051377182e-07 wa2=-5.161821280e-06 pa2=8.716767595e-13 b0=0.0 b1=0.0 keta=5.292491321e-02 lketa=-2.127372133e-08 wketa=-2.173885329e-07 pketa=3.671040154e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.361753037e+00 lpclm=3.540264066e-07 wpclm=3.617668951e-06 ppclm=-6.109157558e-13 pdiblc1=-1.376095058e+00 lpdiblc1=3.103208367e-07 wpdiblc1=3.171057399e-06 ppdiblc1=-5.354964629e-13 pdiblc2=-3.076068581e-02 lpdiblc2=6.862893847e-09 wpdiblc2=7.012945227e-08 ppdiblc2=-1.184276061e-14 pdiblcb=4.129851026e+00 lpdiblcb=-7.353389020e-07 wpdiblcb=-7.514164664e-06 ppdiblcb=1.268916987e-12 drout=-4.682108439e+00 ldrout=9.062445604e-07 wdrout=9.260588328e-06 pdrout=-1.563835551e-12 pscbe1=7.967858873e+08 lpscbe1=5.427673004e-01 wpscbe1=5.546344493e+00 ppscbe1=-9.366111945e-7 pscbe2=5.411646669e-09 lpscbe2=6.600005278e-16 wpscbe2=6.744308822e-15 ppscbe2=-1.138911431e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.939693167e+00 lbeta0=8.454816830e-07 wbeta0=8.639674263e-06 pbeta0=-1.458981793e-12 agidl=5.060553448e-09 lagidl=-8.004443770e-16 wagidl=-8.179454176e-15 pagidl=1.381264427e-21 bgidl=1.869343746e+09 lbgidl=-1.468060825e+02 wbgidl=-1.500158735e+03 pbgidl=2.533318057e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.166979554e-01 lkt1=2.261084232e-08 wkt1=2.310520930e-07 pkt1=-3.901776694e-14 kt2=-7.305882895e-02 lkt2=4.097939491e-09 wkt2=4.187537479e-08 pkt2=-7.071494540e-15 at=7.516085239e+05 lat=-1.252573176e-01 wat=-1.279959632e+00 pat=2.161467830e-7 ute=4.162836676e-01 lute=-7.367522280e-08 wute=-7.528606936e-07 pute=1.271355853e-13 ua1=2.107320144e-08 lua1=-3.414521237e-15 wua1=-3.489176862e-14 pua1=5.892172967e-21 ub1=-2.173378374e-17 lub1=3.590958692e-24 wub1=3.669471972e-23 pub1=-6.196637320e-30 uc1=-2.013766689e-09 luc1=3.356300865e-16 wuc1=3.429683550e-15 puc1=-5.791706611e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.246317546e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.998280012e-08 wvth0=3.495045746e-07 pvth0=-6.496241528e-14 k1=4.071238096e-01 lk1=1.030285673e-07 wk1=-1.856282002e-07 pk1=3.450271357e-14 k2=1.863348031e-01 lk2=-6.227188854e-08 wk2=-3.889440320e-08 pk2=7.229302723e-15 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.081497471e+00 ldsub=-2.823726010e-07 wdsub=-2.328098911e-07 pdsub=4.327237445e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.455985969e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.297067068e-08 wvoff=-1.600085568e-07 pvoff=2.974079045e-14 nfactor='9.066182867e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.067839097e-06 wnfactor=-2.934364304e-07 pnfactor=5.454102932e-14 eta0=-5.351278317e-03 leta0=9.207094210e-08 weta0=3.883159789e-06 peta0=-7.217629099e-13 etab=-1.261599351e+00 letab=2.343773026e-07 wetab=2.577547717e-06 petab=-4.790887941e-13 u0=1.676608934e-02 lu0=-2.353214383e-09 wu0=-1.783503571e-08 pu0=3.314998087e-15 ua=4.099998028e-09 lua=-1.119298659e-15 wua=-9.748913973e-15 pua=1.812030640e-21 ub=-1.495708114e-18 lub=6.042397150e-25 wub=5.376526352e-24 pub=-9.993349530e-31 uc=-5.736685821e-11 luc=9.115493085e-18 wuc=1.160732617e-16 puc=-2.157453716e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.168656581e+05 lvsat=-9.993123173e-02 wvsat=-8.232037424e-01 pvsat=1.530088796e-7 a0=-6.898956592e+00 la0=1.423217109e-06 wa0=1.415145174e-05 pa0=-2.630330335e-12 ags=1.249999831e+00 lags=2.634467666e-14 a1=0.0 a2=-1.595100384e+00 la2=4.196897862e-07 wa2=3.575474744e-06 pa2=-6.645734907e-13 b0=5.904230970e-23 lb0=-1.097419410e-29 wb0=-1.207782477e-28 pb0=2.244905289e-35 b1=0.0 keta=-5.965750302e-01 lketa=9.730722563e-08 wketa=4.075606500e-07 pketa=-7.575329802e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.349047126e+00 lpclm=-3.000604809e-07 wpclm=-2.175207151e-06 ppclm=4.043057532e-13 pdiblc1=2.189823244e+00 lpdiblc1=-3.212366621e-07 wpdiblc1=-3.333371279e-07 ppdiblc1=6.195737197e-14 pdiblc2=5.719952706e-02 lpdiblc2=-8.795389203e-09 wpdiblc2=-2.902534233e-08 ppdiblc2=5.394940379e-15 pdiblcb=3.433942151e+01 lpdiblcb=-6.424417713e-06 wpdiblcb=-6.098588770e-05 ppdiblcb=1.133544695e-11 drout=-9.552668171e-01 ldrout=3.047673812e-07 wdrout=-3.311541533e-12 pdrout=6.155162247e-19 pscbe1=7.895341633e+08 lpscbe1=1.945285156e+00 wpscbe1=2.140915229e+01 ppscbe1=-3.979319137e-6 pscbe2=-3.358980641e-08 lpscbe2=7.975642307e-15 wpscbe2=8.798849792e-14 ppscbe2=-1.635442211e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.969833793e+01 lbeta0=-1.998463693e-06 wbeta0=-1.235519942e-05 pbeta0=2.296460916e-12 agidl=1.642108846e-08 lagidl=-2.992607077e-15 wagidl=-3.092114238e-14 pagidl=5.747312734e-21 bgidl=9.999998475e+08 lbgidl=2.376335716e-5 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.000699791e+00 lkt1=1.211481478e-06 wkt1=1.453792164e-05 pkt1=-2.702163496e-12 kt2=-2.619595634e-02 lkt2=-4.199926541e-09 wkt2=-1.487305687e-13 pkt2=2.764455076e-20 at=1.811172815e+05 lat=-3.182965858e-02 wat=-4.694036583e-01 pat=8.724805796e-8 ute=1.325677166e+00 lute=-2.501210147e-07 wute=8.724083407e-13 pute=-1.621545381e-19 ua1=4.796705996e-09 lua1=-7.329459926e-16 wua1=-3.438854770e-15 pua1=6.391799362e-22 ub1=-2.170212456e-18 lub1=3.161764694e-25 wub1=1.522202020e-30 pub1=-2.829316898e-37 uc1=-7.606959999e-10 luc1=1.365094343e-16 wuc1=1.501632464e-15 puc1=-2.791084260e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos lmin=2.0e-05 lmax=0.0001 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.100659040e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.397772846e-7 k1=4.212606180e-01 lk1=1.291674424e-6 k2=3.716651602e-02 lk2=-5.420869610e-7 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.302605061e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.880721963e-7 nfactor='7.461046316e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.114104823e-5 eta0=0.08 etab=-0.07 u0=1.445963384e-02 lu0=-2.837462552e-8 ua=-6.324241445e-10 lua=4.503683210e-16 ub=1.868978521e-18 lub=-4.055915651e-24 uc=-7.214960068e-11 luc=-7.406433888e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160312.5 a0=1.684311541e+00 la0=-1.357442978e-6 ags=5.136952411e-01 lags=-7.041817269e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-5.480298045e-02 lketa=4.710778082e-07 wketa=8.881784197e-22 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.042722157e-01 lpclm=-2.880916892e-6 pdiblc1=0.39 pdiblc2=1.362535913e-04 lpdiblc2=3.013041483e-9 pdiblcb=-3.448804924e-03 lpdiblcb=3.834829377e-8 drout=0.56 pscbe1=7.008738872e+08 lpscbe1=1.786719392e+3 pscbe2=9.665980000e-09 lpscbe2=-6.105490408e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=5.681322036e-10 lalpha0=-9.357433760e-15 alpha1=-2.464203913e-11 lalpha1=2.491453517e-15 walpha1=1.227846222e-31 palpha1=2.584939414e-35 beta0=3.268447993e+00 lbeta0=-5.365972042e-06 wbeta0=-5.684341886e-20 agidl=5.811380381e-09 lagidl=-1.111856617e-13 bgidl=1.562948962e+09 lbgidl=-1.125271361e+4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.257308181e-01 lkt1=-5.958518612e-7 kt2=-0.037961 at=0.0 ute=-3.559870728e-01 lute=5.256487698e-7 ua1=2.139764998e-09 lua1=7.182700633e-15 ub1=-7.306057684e-19 lub1=-1.899330897e-23 uc1=4.338507642e-11 luc1=7.645641303e-15 puc1=5.293955920e-35 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0886635+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.4858803 k2=0.010047076 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.64967492+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='8.0184089+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0130401126 ua=-6.0989319e-10 ub=1.66606982e-18 uc=-1.0920239e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160312.5 a0=1.6164016 ags=0.47846655 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-0.031235975 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.060146165 pdiblc1=0.39 pdiblc2=0.00028698955 pdiblcb=-0.0015303226 drout=0.56 pscbe1=790259600.0 pscbe2=9.3605355e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.0 agidl=2.4900183e-10 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.45554 kt2=-0.037961 at=0.0 ute=-0.32969 ua1=2.4991e-9 ub1=-1.6808e-18 uc1=4.2588e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.093883435e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.170138215e-8 k1=4.522972755e-01 lk1=2.682904169e-7 k2=2.243897693e-02 lk2=-9.899728555e-08 pk2=8.881784197e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.724699858e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.821068169e-7 nfactor='8.375619887e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.853712138e-6 eta0=0.08 etab=-0.07 u0=1.610008706e-02 lu0=-2.444573819e-8 ua=-1.211989359e-10 lua=-3.904114865e-15 ub=1.642518584e-18 lub=1.881477614e-25 uc=-1.423307551e-10 luc=2.646582022e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.212579461e+05 lvsat=-4.868852462e-1 a0=1.673710294e+00 la0=-4.578317032e-7 ags=4.558541944e-01 lags=1.806471690e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-3.743565127e-02 lketa=4.952840774e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.109267259e-01 lpclm=4.562227086e-06 wpclm=-3.552713679e-21 ppclm=2.131628207e-26 pdiblc1=0.39 pdiblc2=3.587787891e-04 lpdiblc2=-5.735148984e-10 pdiblcb=-4.459427061e-04 lpdiblcb=-8.662970003e-9 drout=0.56 pscbe1=7.805463027e+08 lpscbe1=7.759826970e+1 pscbe2=9.153007757e-09 lpscbe2=1.657912159e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-6.819567689e-01 lbeta0=2.941467397e-5 agidl=-4.042535850e-10 lagidl=5.218772587e-15 pagidl=-2.646977960e-35 bgidl=8.022575536e+08 lbgidl=1.579738698e+3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.101376581e-01 lkt1=4.361735931e-7 kt2=-3.138933667e-02 lkt2=-5.250016399e-8 at=-1.789107917e+05 lat=1.429295056e+0 ute=1.617288118e-01 lute=-3.925881003e-6 ua1=5.328096354e-09 lua1=-2.260048410e-14 ub1=-4.224512371e-18 lub1=2.032138745e-23 uc1=7.901037197e-10 luc1=-2.909735948e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.091149793e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.079724093e-8 k1=5.977558582e-01 lk1=-3.119249599e-7 k2=-2.975396524e-02 lk2=1.091935757e-07 wk2=-2.220446049e-22 pk2=5.551115123e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.915414784e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.581805218e-7 nfactor='8.421149226e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.035322754e-6 eta0=0.08 etab=-0.07 u0=8.149894523e-03 lu0=7.266546324e-9 ua=-1.665485757e-09 lua=2.255844507e-15 ub=2.098150966e-18 lub=-1.629310578e-24 uc=-6.694967090e-11 luc=-3.602714318e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.447013512e+05 lvsat=-1.815109412e-1 a0=1.964587897e+00 la0=-1.618104650e-6 ags=6.476342087e-01 lags=-5.843383766e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-4.118284482e-02 lketa=6.447547569e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.336218480e-01 lpclm=-1.199889384e-6 pdiblc1=0.39 pdiblc2=0.000215 pdiblcb=1.963998626e-02 lpdiblcb=-8.878312947e-08 wpdiblcb=-1.110223025e-22 ppdiblcb=-6.661338148e-28 drout=0.56 pscbe1=800000000.0 pscbe2=1.671893803e-08 lpscbe2=-2.852160011e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.565947440e+00 lbeta0=4.492596311e-6 agidl=5.125510518e-10 lagidl=1.561758076e-15 bgidl=1.143013757e+09 lbgidl=2.205064997e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.434839429e-01 lkt1=-2.285864121e-7 kt2=-4.017360155e-02 lkt2=-1.746087337e-8 at=2.745973838e+05 lat=-3.796900997e-1 ute=-1.640382899e+00 lute=3.262508336e-6 ua1=-3.274541222e-09 lua1=1.171431885e-14 wua1=2.646977960e-29 pua1=2.646977960e-35 ub1=3.170152177e-18 lub1=-9.174968124e-24 wub1=2.465190329e-38 pub1=-9.860761315e-44 uc1=9.216446460e-11 luc1=-1.257469911e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.090845143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.019133174e-8 k1=4.322967437e-01 lk1=1.715170913e-8 k2=2.844424485e-02 lk2=-6.555098444e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.916658762e-01 ldsub=3.347946888e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.722230050e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.087158959e-8 nfactor='8.494631950e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.181470339e-6 eta0=-5.744849986e-02 leta0=2.733671979e-7 etab=6.842919891e-01 letab=-1.500188708e-06 wetab=5.329070518e-21 petab=-1.776356839e-27 u0=1.359424468e-02 lu0=-3.561558378e-9 ua=-1.917591780e-10 lua=-6.752060745e-16 ub=1.151418582e-18 lub=2.536170597e-25 uc=-1.214437714e-10 luc=7.235453841e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.038194939e+04 lvsat=2.596678738e-2 a0=1.099283968e+00 la0=1.028723755e-7 ags=1.353546988e-01 lags=4.345189724e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-2.629453859e-03 lketa=-1.220220699e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.108255342e-02 lpclm=5.752552428e-7 pdiblc1=4.088045794e-01 lpdiblc1=-3.739986375e-8 pdiblc2=2.392950000e-06 lpdiblc2=4.228477835e-10 pdiblcb=-0.025 drout=1.344068365e-01 ldrout=8.464494752e-7 pscbe1=800000000.0 pscbe2=-4.454152232e-09 lpscbe2=1.358892391e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.794355910e+00 lbeta0=2.049451557e-6 agidl=6.445524780e-10 lagidl=1.299224399e-15 bgidl=1.269088568e+09 lbgidl=-3.023991007e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.444605805e-01 lkt1=-2.775700689e-8 kt2=-6.040588351e-02 lkt2=2.277850526e-8 at=6.493100483e+04 lat=3.730907145e-2 ute=0.0 ua1=2.824339679e-09 lua1=-4.155624112e-16 ub1=-1.527062104e-18 lub1=1.671804431e-25 uc1=1.528486051e-10 luc1=-2.464398577e-16 wuc1=8.271806126e-31 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.084139568e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.356038974e-8 k1=3.328536151e-01 lk1=1.154880357e-7 k2=6.118412774e-02 lk2=-3.893058644e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=4.664626476e-01 ldsub=2.608304055e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.014237749e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.974735493e-8 nfactor='5.907109181e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.227466980e-7 eta0=3.582529886e-01 leta0=-1.377075330e-7 etab=-1.646537114e+00 letab=8.046982669e-7 u0=1.169191212e-02 lu0=-1.680398776e-09 wu0=2.220446049e-22 ua=-5.906662208e-10 lua=-2.807388671e-16 ub=1.291920204e-18 lub=1.146792206e-25 uc=-6.422249855e-11 luc=1.577013837e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.500035228e+04 lvsat=1.622387311e-3 a0=1.225620556e+00 la0=-2.205808617e-8 ags=-8.827609932e-02 lags=6.556607597e-7 a1=0.0 a2=6.044617774e-01 la2=1.933618822e-7 b0=0.0 b1=0.0 keta=1.631183582e-02 lketa=-3.093268012e-08 pketa=2.220446049e-28 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.378830106e-01 lpclm=8.398417474e-8 pdiblc1=-2.440305587e-01 lpdiblc1=6.081692192e-7 pdiblc2=-1.444786656e-04 lpdiblc2=5.680847180e-10 pdiblcb=-4.911716338e-02 lpdiblcb=2.384873935e-8 drout=1.009114736e+00 ldrout=-1.852292549e-8 pscbe1=8.085510012e+08 lpscbe1=-8.455828520e+0 pscbe2=9.336779542e-09 lpscbe2=-4.851479500e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.461134792e+00 lbeta0=4.012239235e-7 agidl=2.424195336e-09 lagidl=-4.606110339e-16 bgidl=1.280411890e+09 lbgidl=-4.143720287e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.540604914e-01 lkt1=-1.826394297e-8 kt2=-2.736871980e-02 lkt2=-9.890954821e-9 at=1.688138884e+05 lat=-6.541759562e-2 ute=1.955480000e-02 lute=-1.933715508e-8 ua1=2.651272672e-09 lua1=-2.444216402e-16 ub1=-1.049425256e-18 lub1=-3.051403071e-25 uc1=-1.219162794e-10 luc1=2.526689368e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.376634204e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.804740468e-8 k1=1.942152608e-01 lk1=1.832641680e-7 k2=1.059965720e-01 lk2=-6.083804605e-08 pk2=-4.440892099e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.418210343e+00 ldsub=-2.044504902e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.252626366e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.140145927e-8 nfactor='5.887005239e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.129184837e-7 eta0=-3.184587778e-01 leta0=1.931165483e-07 weta0=-1.776356839e-21 etab=-3.801533128e-04 letab=-5.848652817e-11 u0=1.221893396e-02 lu0=-1.938043943e-9 ua=-4.416108828e-10 lua=-3.536075502e-16 ub=1.308016311e-18 lub=1.068103164e-25 uc=-5.455131315e-11 luc=1.104218596e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.789834292e+04 lvsat=5.094346627e-3 a0=1.584094753e+00 la0=-1.973053668e-7 ags=1.255670918e+00 lags=-1.354618715e-9 a1=0.0 a2=1.322097146e+00 la2=-1.574685206e-7 b0=0.0 b1=0.0 keta=-2.203352684e-02 lketa=-1.218678267e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.857741658e-01 lpclm=1.168462571e-8 pdiblc1=1.514491131e+00 lpdiblc1=-2.515192790e-07 wpdiblc1=-2.842170943e-20 pdiblc2=-7.449769845e-03 lpdiblc2=4.139422417e-09 wpdiblc2=-2.775557562e-23 ppdiblc2=-2.081668171e-29 pdiblcb=2.139637357e-01 lpdiblcb=-1.047636198e-07 wpdiblcb=-2.359223927e-22 ppdiblcb=-4.475586568e-28 drout=1.245268568e+00 ldrout=-1.339714492e-7 pscbe1=7.828979972e+08 lpscbe1=4.085155538e+0 pscbe2=9.158770415e-09 lpscbe2=3.850852687e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=9.602374377e+00 lbeta0=-1.566938724e-7 agidl=2.591742216e-09 lagidl=-5.425196773e-16 bgidl=1.382591054e+09 lbgidl=-9.138953103e+1 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.996533779e-01 lkt1=4.025051457e-9 kt2=-4.646302380e-02 lkt2=-5.563224232e-10 at=5.901083391e+04 lat=-1.173817637e-2 ute=-2.000000080e-02 lute=3.899890411e-16 ua1=3.391436548e-09 lua1=-6.062655543e-16 ub1=-2.824427839e-18 lub1=5.626052055e-25 uc1=-1.122454153e-10 luc1=2.053909835e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.13880799562893+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.961428255393082 k2=-0.148694456831761 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.562303405039308 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.368212947389937+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='3.3210970722327+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.49 etab=-0.000625 u0=0.0041055503490566 ua=-1.92194558459119e-9 ub=1.75516461966667e-18 uc=-8.324553995283e-12 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=79225.201156122 a0=0.758099999261006 ags=1.24999997272013 a1=0.0 a2=0.662874470440252 b0=0.0 b1=0.0 keta=-0.0730519999606918 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.734690420259434 pdiblc1=0.461536473183962 pdiblc2=0.00987941513820755 pdiblcb=-0.224616327814465 drout=0.684413503600629 pscbe1=800000000.518868 pscbe2=9.31998164677673e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.94639467130503 agidl=3.20550031084906e-10 bgidl=999999975.393082 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.482802992940252 kt2=-0.0487919994941038 at=9870.39612421382 ute=-0.0199999991650943 ua1=8.53380055896226e-10 ub1=-4.69150049528303e-19 uc1=-2.62609955581761e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.65e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.043780707e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.766272205e-08 wvth0=2.550245426e-12 pvth0=-4.740141009e-19 k1=2.995547351e-01 lk1=1.230224312e-07 wk1=-4.638744258e-12 pk1=8.622033931e-19 k2=1.637940389e-01 lk2=-5.808223670e-08 wk2=2.435342125e-12 pk2=-4.526570372e-19 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.946566500e+00 ldsub=-2.572929815e-07 wdsub=2.996034488e-11 pdsub=-5.568729293e-18 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.383262249e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.020595489e-08 wvoff=4.278073220e-12 pvoff=-7.951654695e-19 nfactor='8.896182395e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.036241109e-06 wnfactor=-7.987474896e-11 pnfactor=1.484631957e-17 eta0=2.244936646e+00 leta0=-3.261900743e-07 weta0=1.344066141e-11 peta0=-2.498215743e-18 etab=2.320943525e-01 letab=-4.325554605e-08 wetab=-2.999119890e-12 petab=5.574464145e-19 u0=6.430645205e-03 lu0=-4.321653808e-10 wu0=3.407776283e-14 pu0=-6.334033797e-21 ua=-1.549498325e-09 lua=-6.922677217e-17 wua=-1.877841360e-20 pua=3.490343731e-27 ub=1.620010242e-18 lub=2.512114415e-26 wub=-2.578973141e-29 pub=4.793537375e-36 uc=9.897706192e-12 luc=-3.386971501e-18 wuc=4.957926535e-23 puc=-9.215298052e-30 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.398185148e+05 lvsat=-1.126247921e-02 wvsat=-6.968776360e-07 pvsat=1.295286464e-13 a0=1.301824142e+00 la0=-1.010620064e-07 wa0=4.089757397e-12 pa0=-7.601632177e-19 ags=1.249999831e+00 lags=2.634469354e-14 a1=0.0 a2=4.768820509e-01 la2=3.457041102e-08 wa2=1.627072265e-11 pa2=-3.024239220e-18 b0=-1.094875900e-23 lb0=2.035045836e-30 wb0=-1.196924258e-34 pb0=2.224723122e-41 b1=0.0 keta=-3.603916731e-01 lketa=5.340782504e-08 wketa=-2.547054891e-12 pketa=4.734210934e-19 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.088513738e+00 lpclm=-6.576514013e-08 wpclm=-3.005929216e-12 ppclm=5.587120597e-19 pdiblc1=1.996662586e+00 lpdiblc1=-2.853338906e-07 wpdiblc1=-1.484718064e-11 ppdiblc1=2.759645469e-18 pdiblc2=4.037920184e-02 lpdiblc2=-5.668995354e-09 wpdiblc2=1.809217531e-13 ppdiblc2=-3.362792622e-20 pdiblcb=-1.001973283e+00 lpdiblcb=1.444873373e-07 wpdiblcb=6.702776716e-13 ppdiblcb=-1.245845063e-19 drout=-9.552857037e-01 ldrout=3.047708917e-07 wdrout=2.927942791e-11 pdrout=-5.442167264e-18 pscbe1=8.019400484e+08 lpscbe1=-3.605966932e-01 wpscbe1=1.284166687e-03 ppscbe1=-2.386880646e-10 pscbe2=1.739956503e-08 lpscbe2=-1.501752163e-15 wpscbe2=1.167985276e-19 ppscbe2=-2.170934231e-26 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.253849864e+01 lbeta0=-6.676643648e-07 wbeta0=-2.323415902e-11 pbeta0=4.318533342e-18 agidl=-1.497745042e-09 lagidl=3.379665052e-16 wagidl=-9.082793639e-21 pagidl=1.688218853e-27 bgidl=9.999998475e+08 lbgidl=2.376335144e-5 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.424046556e+00 lkt1=-3.544261257e-07 wkt1=-5.998452821e-12 pkt1=1.114932431e-18 kt2=-2.619680459e-02 lkt2=-4.199768877e-09 wkt2=1.315020793e-12 pkt2=-2.444229148e-19 at=-9.090145530e+04 lat=1.873046402e-02 wat=-2.141696499e-06 pat=3.980771280e-13 ute=1.325682142e+00 lute=-2.501219395e-07 wute=-7.713512574e-12 pute=1.433710575e-18 ua1=2.803882499e-09 lua1=-3.625398891e-16 wua1=5.298384738e-21 pua1=-9.848107706e-28 ub1=-2.170203774e-18 lub1=3.161748558e-25 wub1=-1.345874841e-29 pub1=2.501577567e-36 uc1=1.095003338e-10 luc1=-2.523395829e-17 wuc1=2.525776211e-21 puc1=-4.694660250e-28 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos lmin=2.0e-05 lmax=0.0001 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.118298027e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.209164525e-06 wvth0=2.990905505e-08 pvth0=2.456857609e-12 k1=1.728409333e-01 lk1=8.824441367e-06 wk1=4.212258826e-07 pk1=-1.277272535e-11 k2=1.375340493e-01 lk2=-3.314597553e-06 wk2=-1.701853975e-07 pk2=4.701129955e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.040447419e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.190209519e-06 wvoff=-4.445202643e-08 pvoff=-4.371791199e-12 nfactor='5.906875958e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.726799619e-05 wnfactor=2.635285452e-06 pnfactor=-1.038898776e-11 eta0=0.08 etab=-0.07 u0=1.630851505e-02 lu0=1.669338648e-07 wu0=-3.135003647e-09 pu0=-3.311693730e-13 ua=-7.471786972e-10 lua=5.890308438e-15 wua=1.945803441e-16 pua=-9.224082141e-21 ub=2.011695620e-18 lub=3.601695043e-23 wub=-2.419942532e-25 pub=-6.794843333e-29 uc=8.319917263e-11 luc=-6.350317454e-15 wuc=-2.634127977e-16 puc=9.511886758e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.603104088e+05 lvsat=2.090945812e-04 wvsat=3.545848372e-06 pvsat=-3.545453719e-10 a0=1.685114900e+00 la0=1.674986338e-05 wa0=-1.362194143e-09 pa0=-3.070314703e-11 ags=3.582735617e-01 lags=2.427120081e-05 wags=2.635364189e-07 pags=-4.234880809e-11 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-1.091357611e-01 lketa=-4.079618329e-07 wketa=9.212785820e-08 pketa=1.490518954e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=7.543676277e-01 lpclm=-1.928451140e-05 wpclm=-9.327538827e-07 ppclm=2.781429574e-11 pdiblc1=0.39 pdiblc2=-3.413474094e-04 lpdiblc2=1.039773684e-08 wpdiblc2=8.098307639e-10 ppdiblc2=-1.252165192e-14 pdiblcb=-1.383443847e-01 lpdiblcb=1.301259714e-05 wpdiblcb=2.287319127e-07 ppdiblcb=-2.199942178e-11 drout=0.56 pscbe1=4.097397702e+08 lpscbe1=6.957618348e+03 wpscbe1=4.936534138e+02 ppscbe1=-8.767890029e-3 pscbe2=7.396955570e-09 lpscbe2=3.025758131e-13 wpscbe2=3.847407743e-15 ppscbe2=-5.234068093e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=2.135321188e-09 lalpha0=-4.068377063e-14 walpha0=-2.657360120e-15 palpha0=5.311762598e-20 alpha1=-4.419122658e-10 lalpha1=1.083221383e-14 walpha1=7.075325764e-16 palpha1=-1.414277669e-20 beta0=6.909590680e+00 lbeta0=-2.975440007e-04 wbeta0=-6.174001644e-06 pbeta0=4.954234933e-10 agidl=1.054526919e-07 lagidl=-8.584492154e-12 wagidl=-1.689539999e-13 pagidl=1.436752490e-17 bgidl=3.447560627e+09 lbgidl=-4.892397119e+04 wbgidl=-3.195589001e+03 pbgidl=6.387621311e-2 cgidl=300.0 egidl=7.570061872e-01 legidl=-6.569330624e-05 wegidl=-1.114034145e-06 pegidl=1.113910153e-10 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.135837395e-01 lkt1=-3.825819494e-06 wkt1=-1.901590537e-07 pkt1=5.476804178e-12 kt2=-5.000407391e-02 lkt2=1.204173351e-06 wkt2=2.042050106e-08 pkt2=-2.041822826e-12 at=0.0 ute=-2.788836306e-01 lute=-1.422671664e-05 wute=-1.307382929e-07 pute=2.501443533e-11 ua1=3.710327627e-10 lua1=8.779917495e-14 wua1=2.999101291e-15 pua1=-1.366950674e-19 ub1=3.257526331e-18 lub1=-1.632812093e-22 wub1=-6.762364526e-24 pub1=2.446577382e-28 uc1=-1.600676817e-09 luc1=6.959378104e-14 wuc1=2.787707516e-15 puc1=-1.050406286e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.178789917e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' wvth0=1.528203356e-7 k1=6.143086784e-01 wk1=-2.177659839e-7 k2=-2.828810839e-02 wk2=6.500198203e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.944732894e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' wvoff=-2.631632992e-7 nfactor='6.770756517e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=2.115546829e-6 eta0=0.08 etab=-0.07 u0=2.465985581e-02 wu0=-1.970269222e-8 ua=-4.524992862e-10 wua=-2.668805660e-16 ub=3.813545872e-18 wub=-3.641307637e-24 uc=-2.344934960e-10 wuc=2.124463558e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.603208694e+05 wvsat=-1.419129094e-5 a0=2.523074394e+00 wa0=-1.537374336e-6 ags=1.572509325e+00 wags=-1.855082997e-6 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-1.295452106e-01 wketa=1.666953027e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-2.103948328e-01 wpclm=4.587352678e-7 pdiblc1=0.39 pdiblc2=1.788289110e-04 wpdiblc2=1.833995591e-10 pdiblcb=5.126477496e-01 wpdiblcb=-8.718516511e-7 drout=0.56 pscbe1=7.578143911e+08 wpscbe1=5.501480994e+1 pscbe2=2.253417009e-08 wpscbe2=-2.233750462e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-7.975893126e+00 wbeta0=1.861096585e-5 agidl=-3.240109123e-07 wagidl=5.498222441e-13 bgidl=1000000000.0 cgidl=300.0 egidl=-2.529488059e+00 wegidl=4.458617801e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.049812269e-01 wkt1=8.383363211e-8 kt2=1.023811843e-02 wkt2=-8.172748559e-8 at=0.0 ute=-9.906155412e-01 wute=1.120679888e-6 ua1=4.763435883e-09 wua1=-3.839457738e-15 ub1=-4.911079965e-18 wub1=5.477333775e-24 uc1=1.880949760e-09 wuc1=-2.467248297e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.182522580e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.981975812e-08 wvth0=1.502984842e-07 pvth0=2.014674311e-14 k1=4.412317095e-01 lk1=1.382689405e-06 wk1=1.876301716e-08 pk1=-1.889599441e-12 k2=3.434970078e-02 lk2=-5.004053146e-07 wk2=-2.019608540e-08 pk2=6.806362850e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.672212293e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.177131657e-07 wvoff=-3.480243069e-07 pvoff=6.779435586e-13 nfactor='5.561537399e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.660294335e-06 wnfactor=4.771620177e-06 pnfactor=-2.121902468e-11 eta0=0.08 etab=-0.07 u0=3.908690492e-02 lu0=-1.152558199e-07 wu0=-3.897695407e-08 pu0=1.539795723e-13 ua=1.800356156e-09 lua=-1.799776925e-14 wua=-3.258231087e-15 pua=2.389751044e-20 ub=3.684350605e-18 lub=1.032124187e-24 wub=-3.462175295e-24 pub=-1.431064994e-30 uc=-3.816433969e-10 luc=1.175561429e-15 wuc=4.057837803e-16 puc=-1.544547551e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.851127815e+04 lvsat=7.334548890e-01 wvsat=2.590006106e-01 pvsat=-2.069235581e-6 a0=2.512905332e+00 la0=8.123931291e-08 wa0=-1.422957570e-06 pa0=-9.140606745e-13 ags=1.556131661e+00 lags=1.308390276e-07 wags=-1.865654678e-06 pags=8.445578024e-14 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-1.599307534e-01 lketa=2.427461510e-07 wketa=2.077053900e-07 pketa=-3.276242562e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-3.024352626e+00 lpclm=2.248034299e-05 wpclm=4.261820251e-06 ppclm=-3.038235153e-11 pdiblc1=0.39 pdiblc2=6.189427901e-03 lpdiblc2=-4.801789395e-08 wpdiblc2=-9.886576909e-09 ppdiblc2=8.044773290e-14 pdiblcb=8.302761565e-01 lpdiblcb=-2.537492052e-06 wpdiblcb=-1.408590667e-06 ppdiblcb=4.287938225e-12 drout=0.56 pscbe1=-7.024619961e+08 lpscbe1=1.166595822e+04 wpscbe1=2.514621498e+03 ppscbe1=-1.964947808e-2 pscbe2=9.644516451e-08 lpscbe2=-5.904653260e-13 wpscbe2=-1.480145014e-13 ppscbe2=1.004017189e-18 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-1.452847448e+01 lbeta0=5.234772057e-05 wbeta0=2.347846005e-05 pbeta0=-3.888577834e-11 agidl=-6.476107460e-07 lagidl=2.585197004e-12 wagidl=1.097417567e-12 pagidl=-4.374667848e-18 bgidl=1.402655322e+08 lbgidl=6.868306898e+03 wbgidl=1.122488235e+03 pbgidl=-8.967412588e-3 cgidl=300.0 egidl=-5.151659567e+00 legidl=2.094818730e-05 wegidl=8.904829498e-06 pegidl=-3.552020724e-11 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-8.573955395e-01 lkt1=2.815392129e-06 wkt1=5.888181033e-07 pkt1=-4.034255293e-12 kt2=2.564819125e-02 lkt2=-1.231090685e-07 wkt2=-9.671408718e-08 pkt2=1.197260119e-13 at=-4.751433594e+05 lat=3.795858529e+00 wat=5.022984589e-01 pat=-4.012797089e-6 ute=1.253668267e+00 lute=-1.792929159e-05 wute=-1.851516563e-06 pute=2.374449106e-11 ua1=2.121980371e-08 lua1=-1.314677833e-13 wua1=-2.694632861e-14 pua1=1.845977875e-19 ub1=-2.108101345e-17 lub1=1.291794966e-22 wub1=2.858225408e-23 pub1=-1.845822047e-28 uc1=3.474085516e-09 luc1=-1.272735444e-14 wuc1=-4.551018581e-15 puc1=1.664696991e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.198597591e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=9.394088729e-08 wvth0=1.821908495e-07 pvth0=-1.070677559e-13 k1=1.116679585e+00 lk1=-1.311584361e-06 wk1=-8.798984869e-07 pk1=1.695044473e-12 k2=-2.021138318e-01 lk2=4.428169765e-07 wk2=2.922571816e-07 pk2=-5.656991782e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.344110573e-01 ldsub=3.966576434e-06 wdsub=1.686145266e-06 pdsub=-6.725814266e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.196706563e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.903877804e-07 wvoff=-1.218657470e-07 pvoff=-2.241735362e-13 nfactor='9.593284507e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.421820752e-06 wnfactor=-1.987498369e-06 pnfactor=5.742220508e-12 eta0=-1.846649205e-01 leta0=1.055713961e-06 weta0=4.487716618e-07 peta0=-1.790091818e-12 etab=1.613778929e-01 letab=-9.229363358e-07 wetab=-3.923294456e-07 petab=1.564951156e-12 u0=5.637639653e-03 lu0=1.816895088e-08 wu0=4.259834627e-09 pu0=-1.848635702e-14 ua=-4.699980971e-09 lua=7.931230499e-15 wua=5.145356843e-15 pua=-9.623309348e-21 ub=5.742820689e-18 lub=-7.178845374e-24 wub=-6.179982164e-24 pub=9.409913290e-30 uc=-3.814362266e-11 luc=-1.946145158e-16 wuc=-4.884416912e-17 puc=2.689042380e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.502281180e+05 lvsat=-7.891639620e-01 wvsat=-5.180579075e-01 pvsat=1.030349830e-6 a0=4.387409540e+00 la0=-7.395914285e-06 wa0=-4.108189679e-06 pa0=9.796981129e-12 ags=2.574502579e+00 lags=-3.931310178e-06 wags=-3.267240400e-06 pags=5.675199020e-12 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-2.005320765e-01 lketa=4.046995508e-07 wketa=2.701960629e-07 pketa=-5.768914267e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.886142155e+00 lpclm=-1.306246232e-05 wpclm=-8.397602387e-06 ppclm=2.011443965e-11 pdiblc1=0.39 pdiblc2=-1.116257839e-02 lpdiblc2=2.119700338e-08 wpdiblc2=1.929207222e-08 ppdiblc2=-3.594210526e-14 pdiblcb=4.120466754e-01 lpdiblcb=-8.692290214e-07 wpdiblcb=-6.653734151e-07 ppdiblcb=1.323341224e-12 drout=0.56 pscbe1=3.610583925e+09 lpscbe1=-5.538221261e+03 wpscbe1=-4.765687936e+03 ppscbe1=9.390729811e-3 pscbe2=-8.202937486e-08 lpscbe2=1.214464098e-13 wpscbe2=1.674398118e-13 ppscbe2=-2.542890569e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-1.407591857e+01 lbeta0=5.054253387e-05 wbeta0=3.330518012e-05 pbeta0=-7.808328723e-11 agidl=-2.391713993e-09 lagidl=1.150216340e-14 wagidl=4.924535704e-15 pagidl=-1.685516996e-20 bgidl=1.621787880e+09 lbgidl=9.587068515e+02 wbgidl=-8.118199350e+02 pbgidl=-1.251708757e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=1.185754887e-01 lkt1=-1.077629426e-06 wkt1=-7.834781375e-07 pkt1=1.439656013e-12 kt2=2.693027371e-02 lkt2=-1.282231287e-07 wkt2=-1.137828072e-07 pkt2=1.878109170e-13 at=8.520883640e+05 lat=-1.498296275e+00 wat=-9.792064107e-01 pat=1.896733240e-6 ute=-6.689477486e+00 lute=1.375488421e-05 wute=8.561355863e-06 pute=-1.779110337e-11 ua1=-2.534903998e-08 lua1=5.428928029e-14 wua1=3.743000574e-14 pua1=-7.219104127e-20 ub1=2.326426416e-17 lub1=-4.770805098e-23 wub1=-3.407201836e-23 pub1=6.533754302e-29 uc1=3.412091491e-10 luc1=-2.307178918e-16 wuc1=-4.222856460e-16 puc1=1.779909686e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.152166987e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.596451615e-09 wvth0=1.039786668e-07 pvth0=4.848610783e-14 k1=6.850095563e-01 lk1=-4.530487916e-07 wk1=-4.285054047e-07 pk1=7.972823134e-13 k2=-6.581041321e-02 lk2=1.717271965e-07 wk2=1.598202718e-07 pk2=-3.022993814e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.534590227e+00 ldsub=-1.938381150e-06 wdsub=-3.633589673e-06 pdsub=3.854446962e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.350466824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.756923027e-07 wvoff=-4.021613905e-07 pvoff=3.332980602e-13 nfactor='8.752044052e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.748702848e-06 wnfactor=-4.364736228e-07 pnfactor=2.657433922e-12 eta0=4.752066603e-01 leta0=-2.566848296e-07 weta0=-9.031818080e-07 peta0=8.987678790e-13 etab=2.443710575e-01 letab=-1.087998951e-06 wetab=7.459396098e-07 petab=-6.989180207e-13 u0=1.584830128e-02 lu0=-2.138727709e-09 wu0=-3.822027955e-09 pu0=-2.412582985e-15 ua=2.013489644e-10 lua=-1.816877568e-15 wua=-6.665628147e-16 pua=1.935843302e-21 ub=1.027159610e-18 lub=2.199991475e-24 wub=2.106962456e-25 pub=-3.300315278e-30 uc=-2.772127238e-10 luc=2.808628473e-16 wuc=2.641252626e-16 puc=-3.535512757e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-2.338136527e+04 lvsat=1.527837310e-01 wvsat=1.081184791e-01 pvsat=-2.150335996e-7 a0=1.636421754e-01 la0=1.004609912e-06 wa0=1.586494808e-06 pa0=-1.529006005e-12 ags=1.789740124e-01 lags=8.330847224e-07 wags=-7.396186791e-08 pags=-6.758168541e-13 a1=0.0 a2=1.462064550e+00 la2=-1.316760322e-06 wa2=-1.122611217e-06 pa2=2.232727770e-12 b0=0.0 b1=0.0 keta=2.488727691e-02 lketa=-4.363023861e-08 wketa=-4.665797406e-08 pketa=5.329006183e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.364808545e+00 lpclm=1.358735996e-06 wpclm=2.383859876e-06 ppclm=-1.328487202e-12 pdiblc1=-6.902237986e-01 lpdiblc1=2.148424706e-06 wpdiblc1=1.863536696e-06 ppdiblc1=-3.706332229e-12 pdiblc2=-1.429128003e-03 lpdiblc2=1.838435909e-09 wpdiblc2=2.427318422e-09 ppdiblc2=-2.400302368e-15 pdiblcb=-0.025 drout=1.662427097e-01 ldrout=7.831320619e-07 wdrout=-5.398160712e-08 pdrout=1.073623989e-13 pscbe1=8.063185820e+08 lpscbe1=3.909795145e+01 wpscbe1=-1.071392670e+01 ppscbe1=-6.629534663e-5 pscbe2=-5.125104139e-08 lpscbe2=6.023230573e-14 wpscbe2=7.934983478e-14 ppscbe2=-7.908954437e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=9.811074221e+00 lbeta0=3.034410532e-06 wbeta0=-5.115213936e-06 pbeta0=-1.670118107e-12 agidl=2.003070137e-09 lagidl=2.761509089e-15 wagidl=-2.303532430e-15 pagidl=-2.479482091e-21 bgidl=2.169929479e+09 lbgidl=-1.314755302e+02 wbgidl=-1.527485666e+03 pbgidl=1.716573447e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.961606329e-01 lkt1=-5.388619587e-08 wkt1=-8.189845366e-08 pkt1=4.430522768e-14 kt2=-7.474559650e-02 lkt2=7.399695926e-08 wkt2=2.431473282e-08 pkt2=-8.684713741e-14 at=-4.051388487e+04 lat=2.769735598e-01 wat=1.787946748e-01 pat=-4.063803790e-7 ute=-3.019537603e+00 lute=6.455850877e-06 wute=5.119994390e-06 pute=-1.094668278e-11 ua1=-7.887599455e-09 lua1=1.956074506e-14 wua1=1.816339966e-14 pua1=-3.387226643e-20 ub1=7.362582748e-18 lub1=-1.608167386e-23 wub1=-1.507347738e-23 pub1=2.755191483e-29 uc1=1.083744252e-09 luc1=-1.707523682e-15 wuc1=-1.578447138e-15 puc1=2.477445876e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.166980640e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.624522896e-08 wvth0=1.404671438e-07 pvth0=1.240374755e-14 k1=-2.814058615e-01 lk1=5.026104226e-07 wk1=1.041551882e-06 pk1=-6.564132359e-13 k2=2.783693339e-01 lk2=-1.686218301e-07 wk2=-3.682640137e-07 pk2=2.199073260e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.255588468e+00 ldsub=2.798482856e-06 wdsub=4.615569756e-06 pdsub=-4.302899323e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.083651404e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.302879152e-09 wvoff=-1.577922679e-07 pvoff=9.164876602e-14 nfactor='2.682214290e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.253569708e-06 wnfactor=5.468202725e-06 pnfactor=-3.181523378e-12 eta0=1.704860769e+00 leta0=-1.472652888e-06 weta0=-2.283337777e-06 peta0=2.263562712e-12 etab=-1.692616665e+00 letab=8.274300984e-07 wetab=7.813350071e-08 petab=-3.854459355e-14 u0=2.401827946e-02 lu0=-1.021777403e-08 wu0=-2.090085964e-08 pu0=1.447616130e-14 ua=2.967851474e-11 lua=-1.647117811e-15 wua=-1.051870181e-15 pua=2.316862197e-21 ub=3.364902026e-18 lub=-1.117318676e-25 wub=-3.514993583e-24 pub=3.839076222e-31 uc=5.203953773e-11 luc=-4.472483652e-17 wuc=-1.971364665e-16 puc=1.025766103e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.150824111e+05 lvsat=1.586105646e-02 wvsat=-8.492024075e-02 pvsat=-2.414340066e-8 a0=-3.401710156e-01 la0=1.502815662e-06 wa0=2.654990636e-06 pa0=-2.585609475e-12 ags=7.856307014e-01 lags=2.331801224e-07 wags=-1.481815597e-06 pags=7.163674632e-13 a1=0.0 a2=-7.520729984e-01 la2=8.727338758e-07 wa2=2.300170210e-06 pa2=-1.151958099e-12 b0=0.0 b1=0.0 keta=3.813442977e-02 lketa=-5.672995066e-08 wketa=-3.700287040e-08 pketa=4.374241947e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-2.907425967e+00 lpclm=2.884184086e-06 wpclm=5.841941700e-06 ppclm=-4.748080575e-12 pdiblc1=-1.283195189e+00 lpdiblc1=2.734796325e-06 wpdiblc1=1.762030408e-06 ppdiblc1=-3.605955706e-12 pdiblc2=-3.343804387e-03 lpdiblc2=3.731801944e-09 wpdiblc2=5.424847079e-09 ppdiblc2=-5.364468531e-15 pdiblcb=-1.119480211e-01 lpdiblcb=8.598028965e-08 wpdiblcb=1.065373847e-07 ppdiblcb=-1.053516236e-13 drout=1.039628582e+00 ldrout=-8.053302554e-08 wdrout=-5.173994838e-08 pdrout=1.051456899e-13 pscbe1=9.278700197e+08 lpscbe1=-8.110061869e+01 wpscbe1=-2.023199528e+02 ppscbe1=1.231781044e-4 pscbe2=1.036804785e-08 lpscbe2=-7.009630481e-16 wpscbe2=-1.748641236e-15 ppscbe2=1.106305612e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.466161651e+01 lbeta0=-1.762145218e-06 wbeta0=-1.051367321e-05 pbeta0=3.668256311e-12 agidl=6.432462976e-09 lagidl=-1.618584607e-15 wagidl=-6.796506792e-15 pagidl=1.963485467e-21 bgidl=2.219160434e+09 lbgidl=-1.801585457e+02 wbgidl=-1.591762685e+03 pbgidl=2.352189607e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.634902094e-01 lkt1=1.115810025e-07 wkt1=1.855514374e-07 pkt1=-2.201679461e-13 kt2=9.559689512e-02 lkt2=-9.444962043e-08 wkt2=-2.085032019e-07 pkt2=1.433795337e-13 at=4.398981526e+05 lat=-1.980914917e-01 wat=-4.596564423e-01 pat=2.249647771e-7 ute=6.374961427e+00 lute=-2.834087378e-06 wute=-1.077636729e-05 pute=4.772752402e-12 ua1=2.277750131e-08 lua1=-1.076305313e-14 wua1=-3.412647606e-14 pua1=1.783562297e-20 ub1=-1.846974694e-17 lub1=9.463142001e-24 wub1=2.953828070e-23 pub1=-1.656331438e-29 uc1=-1.612488626e-09 luc1=9.587001245e-16 wuc1=2.527447264e-15 puc1=-1.582749922e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-7.068487552e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.086994456e-07 wvth0=-3.913744243e-07 pvth0=2.724051350e-13 k1=-8.181497841e-01 lk1=7.650084241e-07 wk1=1.716588442e-06 pk1=-9.864183589e-13 k2=5.198290321e-01 lk2=-2.866642327e-07 wk2=-7.017034236e-07 pk2=3.829158503e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=7.051200765e+00 ldsub=-1.751327196e-06 wdsub=-9.551422486e-06 pdsub=2.622918174e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.656506321e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.258927915e-08 wvoff=6.848277356e-08 pvoff=-1.897031352e-14 nfactor='6.314762081e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.222739302e-07 wnfactor=-7.253139129e-07 pnfactor=-1.536988991e-13 eta0=-3.024975615e+00 leta0=8.396222251e-07 weta0=4.589229492e-06 peta0=-1.096229249e-12 etab=2.418731793e-03 letab=-1.221856194e-09 wetab=-4.745851160e-09 petab=1.972635199e-15 u0=1.564970892e-02 lu0=-6.126630953e-09 wu0=-5.817297505e-09 pu0=7.102260283e-15 ua=-1.685710765e-09 lua=-8.085154534e-16 wua=2.109523131e-15 pua=7.713518487e-22 ub=4.199311452e-18 lub=-5.196496039e-25 wub=-4.902543649e-24 pub=1.062239223e-30 uc=-4.240296082e-11 luc=1.445267744e-18 wuc=-2.059901347e-17 puc=1.627274566e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.831892051e+05 lvsat=-1.743431192e-02 wvsat=-2.124459423e-01 pvsat=3.820008907e-8 a0=4.093929001e+00 la0=-6.648828128e-07 wa0=-4.255730168e-06 pa0=7.928346043e-13 ags=2.162616775e+00 lags=-4.399870593e-07 wags=-1.537837347e-06 pags=7.437548161e-13 a1=0.0 a2=1.825532881e+00 la2=-3.873803105e-07 wa2=-8.536367079e-07 pa2=3.898434891e-13 b0=0.0 b1=0.0 keta=4.456765088e-02 lketa=-5.987495946e-08 wketa=-1.129304222e-07 pketa=8.086112170e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.841918725e+00 lpclm=-9.042380533e-07 wpclm=-7.047250150e-06 ppclm=1.553058645e-12 pdiblc1=7.820230090e+00 lpdiblc1=-1.715595191e-06 wpdiblc1=-1.069214971e-05 ppdiblc1=2.482519326e-12 pdiblc2=-3.245454199e-03 lpdiblc2=3.683721488e-09 wpdiblc2=-7.128930104e-09 ppdiblc2=7.726965207e-16 pdiblcb=3.656277649e-01 lpdiblcb=-1.474921849e-07 wpdiblcb=-2.571648646e-07 ppdiblcb=7.245149502e-14 drout=4.320364309e-01 ldrout=2.165005493e-07 wdrout=1.378934302e-06 pdrout=-5.942680310e-13 pscbe1=7.255521866e+08 lpscbe1=1.780650037e+01 wpscbe1=9.723681804e+01 ppscbe1=-2.326621417e-5 pscbe2=8.037511926e-09 lpscbe2=4.383660503e-16 wpscbe2=1.901230561e-15 ppscbe2=-6.780072136e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.310671459e+01 lbeta0=-1.002000316e-06 wbeta0=-5.942036353e-06 pbeta0=1.433320203e-12 agidl=1.402101091e-08 lagidl=-5.328398034e-15 wagidl=-1.937971944e-14 pagidl=8.115040631e-21 bgidl=3.496250376e+09 lbgidl=-8.044895054e+02 wbgidl=-3.583967246e+03 pbgidl=1.209148005e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.049450766e-01 lkt1=-1.481395661e-08 wkt1=-3.301516792e-07 pkt1=3.194383654e-14 kt2=-1.576485041e-01 lkt2=2.935445787e-08 wkt2=1.885285464e-07 pkt2=-5.071737710e-14 at=2.573329861e+05 lat=-1.088408588e-01 wat=-3.362794043e-01 pat=1.646494445e-7 ute=-1.551221188e+00 lute=1.040785517e-06 wute=2.596372332e-06 pute=-1.764778819e-12 ua1=-1.127402449e-09 lua1=9.233371685e-16 wua1=7.662242818e-15 pua1=-2.593628028e-21 ub1=3.127765906e-18 lub1=-1.095234105e-24 wub1=-1.009267066e-23 pub1=2.811068807e-30 uc1=4.591558542e-10 luc1=-5.406471267e-17 wuc1=-9.688805635e-16 puc1=1.264998632e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-2.645606438e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.725176734e-07 wvth0=2.554960589e-06 pvth0=-4.620869624e-13 k1=7.210832963e+00 lk1=-1.234922952e-06 wk1=-1.059662811e-05 pk1=2.093962526e-12 k2=-2.543023256e+00 lk2=4.766263424e-07 wk2=4.059876588e-06 pk2=-8.081781119e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.332924860e+00 ldsub=1.036889841e-06 wdsub=8.300456742e-06 pdsub=-1.758173227e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.228934242e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-8.942020987e-08 wvoff=-6.035118949e-07 pvoff=1.516228751e-13 nfactor='-2.054619694e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.108886388e-06 wnfactor=5.979711095e-06 pnfactor=-1.880252155e-12 eta0=-2.416206241e+00 leta0=7.436109908e-07 weta0=4.927827239e-06 peta0=-1.260883156e-12 etab=-2.396507037e-01 letab=6.062949270e-08 wetab=4.052972418e-07 petab=-1.028047017e-13 u0=-5.008474985e-02 lu0=1.025682238e-08 wu0=9.188626520e-08 pu0=-1.739169368e-14 ua=-1.416655940e-08 lua=2.327418522e-15 wua=2.076223657e-14 pua=-3.946422049e-21 ub=3.502293763e-18 lub=-3.782863280e-25 wub=-2.962470612e-24 pub=6.414306201e-31 uc=-1.827144559e-10 luc=3.744962740e-17 wuc=2.956993542e-16 puc=-6.350041211e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.678081377e+04 lvsat=3.760864441e-02 wvsat=1.967023510e-01 pvsat=-6.377004485e-8 a0=1.895212042e+00 la0=-1.496157623e-07 wa0=-1.928112195e-06 pa0=2.536917781e-13 ags=-2.146985229e+00 lags=6.313976225e-07 wags=5.760002842e-06 pags=-1.070611699e-12 a1=0.0 a2=-1.120302326e+00 la2=3.388013000e-07 wa2=3.023593805e-06 pa2=-5.744789379e-13 b0=0.0 b1=0.0 keta=-3.324608183e-01 lketa=3.233410879e-08 wketa=4.398592993e-07 pketa=-5.482642622e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.798236115e+00 lpclm=-1.898041755e-07 wpclm=-1.803371477e-06 ppclm=3.218361356e-13 pdiblc1=4.213889025e-01 lpdiblc1=5.545010798e-08 wpdiblc1=6.807510406e-08 ppdiblc1=-9.402242300e-14 pdiblc2=3.004518231e-04 lpdiblc2=3.038595145e-09 wpdiblc2=1.624230093e-08 ppdiblc2=-5.152308776e-15 pdiblcb=-3.275013682e-01 lpdiblcb=1.936198095e-08 wpdiblcb=1.744541379e-07 ppdiblcb=-3.283060087e-14 drout=2.603263332e+00 ldrout=-3.236432763e-07 wdrout=-3.253643984e-06 pdrout=5.487766594e-13 pscbe1=8.003542628e+08 lpscbe1=-6.584640191e-02 wpscbe1=-6.006948682e-01 ppscbe1=1.116506077e-7 pscbe2=1.055147437e-08 lpscbe2=-1.736837026e-16 wpscbe2=-2.088146159e-15 ppscbe2=2.945019071e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.269033156e+00 lbeta0=1.187986454e-06 wbeta0=7.931037088e-06 pbeta0=-2.014375967e-12 agidl=-3.398710369e-08 lagidl=6.576224589e-15 wagidl=5.817281242e-14 pagidl=-1.115079109e-20 bgidl=-2.186116388e+09 lbgidl=5.922034331e+02 wbgidl=5.402449000e+03 pbgidl=-1.004153170e-3 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.372318797e+00 lkt1=2.572406713e-07 wkt1=1.508282566e-06 pkt1=-4.361829416e-13 kt2=-3.615905713e-02 lkt2=3.580634082e-10 wkt2=-2.142069499e-08 pkt2=-6.071401923e-16 at=-5.786981700e+05 lat=9.732840140e-02 wat=9.979898092e-01 pat=-1.650321786e-7 ute=8.007161163e+00 lute=-1.330846717e-06 wute=-1.361103106e-05 pute=2.256612971e-12 ua1=3.983878706e-09 lua1=-3.187738951e-16 wua1=-5.308142382e-15 pua1=5.405200295e-22 ub1=-1.170777320e-18 lub1=-7.331192822e-26 wub1=1.189694635e-24 pub1=1.243093183e-31 uc1=6.884804967e-10 luc1=-1.165897090e-16 wuc1=-1.211931399e-15 puc1=1.976920756e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.65e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-7.662716023e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.679429258e-08 wvth0=-4.705479937e-07 pvth0=1.002643179e-13 k1=-2.310853057e+00 lk1=5.348728284e-07 wk1=4.426260242e-06 pk1=-6.983417319e-13 k2=1.379903914e+00 lk2=-2.525281308e-07 wk2=-2.062060224e-06 pk2=3.297062832e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=7.264155629e+00 ldsub=-1.118659509e-06 wdsub=-9.016591154e-06 pdsub=1.460546466e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.667753091e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.182808371e-07 wvoff=1.745523120e-06 pvoff=-2.849922631e-13 nfactor='2.999932779e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.505277885e-06 wnfactor=-3.578303748e-05 pnfactor=5.882189923e-12 eta0=9.214556518e+00 leta0=-1.418198883e-06 weta0=-1.181782735e-05 peta0=1.851631662e-12 etab=1.098339872e+00 letab=-1.880628155e-07 wetab=-1.468827959e-06 petab=2.455389493e-13 u0=1.520704066e-02 lu0=-1.878962721e-09 wu0=-1.488141513e-08 pu0=2.453215066e-15 ua=-2.554588734e-11 lua=-3.009716603e-16 wua=-2.584066058e-15 pua=3.929552211e-22 ub=8.793904358e-19 lub=1.092327134e-25 wub=1.255785448e-24 pub=-1.426166337e-31 uc=9.799438381e-11 luc=-1.472572463e-17 wuc=-1.493786151e-16 puc=1.922623004e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.290003334e+05 lvsat=-4.896609741e-02 wvsat=-4.903437505e-01 pvsat=6.393121404e-8 a0=3.454250056e+00 la0=-4.393941580e-07 wa0=-3.649696643e-06 pa0=5.736826794e-13 ags=1.249999265e+00 lags=1.145400343e-13 wags=9.594276591e-13 pags=-1.495459898e-19 a1=0.0 a2=-1.061225533e-01 la2=1.502957057e-07 wa2=9.885717038e-07 pa2=-1.962293799e-13 b0=-4.760275983e-23 lb0=8.847924970e-30 wb0=6.215121049e-29 pb0=-1.155204549e-35 b1=0.0 keta=-1.407787164e+00 lketa=2.322050167e-07 wketa=1.775984291e-06 pketa=-3.031719784e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.315397010e+00 lpclm=-2.859288711e-07 wpclm=-2.080333273e-06 ppclm=3.733150245e-13 pdiblc1=7.394020791e+00 lpdiblc1=-1.240552981e-06 wpdiblc1=-9.151894161e-06 ppdiblc1=1.619693264e-12 pdiblc2=1.492542833e-01 lpdiblc2=-2.464745351e-08 wpdiblc2=-1.846108024e-07 ppdiblc2=3.218025754e-14 pdiblcb=-3.603082878e+00 lpdiblcb=6.281943163e-07 wpdiblcb=4.410499324e-06 ppdiblcb=-8.201843196e-13 drout=-6.266896325e+00 ldrout=1.325053299e-06 wdrout=9.006513105e-06 pdrout=-1.730018739e-12 pscbe1=8.084381355e+08 lpscbe1=-1.568395831e+00 wpscbe1=-1.101701538e+01 ppscbe1=2.047732102e-6 pscbe2=4.474533569e-08 lpscbe2=-6.529296706e-15 wpscbe2=-4.636797355e-14 ppscbe2=8.524793424e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=2.627803013e+01 lbeta0=-2.902825813e-06 wbeta0=-2.329707509e-05 pbeta0=3.789993244e-12 agidl=-6.511842374e-09 lagidl=1.469397768e-15 wagidl=8.502004664e-15 pagidl=-1.918478053e-21 bgidl=9.999993372e+08 lbgidl=1.033171067e-04 wbgidl=8.654204636e-04 pbgidl=-1.348930874e-10 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=8.302150166e+00 lkt1=-1.540952875e-06 wkt1=-1.166266980e-05 pkt1=2.011901974e-12 kt2=6.400896291e-02 lkt2=-1.826016648e-08 wkt2=-1.529535689e-07 pkt2=2.384087508e-14 at=-4.931973912e+05 lat=8.143637166e-02 wat=6.821396978e-01 pat=-1.063251184e-7 ute=6.697734947e+00 lute=-1.087463666e-06 wute=-9.108978634e-06 pute=1.419816486e-12 ua1=1.074914996e-08 lua1=-1.576234863e-15 wua1=-1.347216501e-14 pua1=2.057966915e-21 ub1=-8.960991806e-18 lub1=1.374655238e-24 wub1=1.151459612e-23 pub1=-1.794780121e-30 uc1=6.514783155e-10 luc1=-1.097121136e-16 wuc1=-9.189872634e-16 puc1=1.432425492e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos lmin=2.0e-05 lmax=0.0001 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.071599519e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.970406590e-07 wvth0=-3.106154497e-08 pvth0=6.208851843e-13 k1=1.059737551e+00 lk1=-1.223758322e-05 wk1=-7.367258537e-07 pk1=1.472631731e-11 k2=-8.856083998e-02 lk2=2.199954043e-06 wk2=1.250090640e-07 pk2=-2.498789929e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.106833681e-04 lcit=-2.012546757e-09 wcit=-1.314544205e-10 pcit=2.627625322e-15 voff='3.241497306e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.870681978e-05 wvoff=-5.065276326e-06 pvoff=1.012491500e-10 nfactor='-2.785378583e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.244941691e-04 wnfactor=4.671394822e-05 pnfactor=-9.337590381e-10 eta0=0.08 etab=-0.07 u0=3.610803541e-02 lu0=-5.304813310e-07 wu0=-2.898569303e-08 pu0=5.793912498e-13 ua=1.386374813e-09 lua=-4.084291533e-14 wua=-2.591034058e-15 pua=5.179184294e-20 ub=4.464896017e-18 lub=-6.876760766e-23 wub=-3.444946661e-24 pub=6.886059097e-29 uc=-1.553851903e-10 luc=1.671235065e-15 wuc=4.808819537e-17 puc=-9.612286857e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.944361679e+05 lvsat=-1.667323953e+01 wvsat=-1.089049396e+00 pvsat=2.176886680e-5 a0=3.269990197e+00 la0=-3.846696516e-05 wa0=-2.070610249e-06 pa0=4.138915909e-11 ags=4.360214229e+00 lags=-8.412410345e-05 wags=-4.961485359e-06 pags=9.917448585e-11 a1=0.0 a2=-9.690507613e-01 la2=3.536132569e-05 wa2=2.309711593e-06 pa2=-4.616852477e-11 b0=1.064552311e-06 lb0=-2.127919775e-11 wb0=-1.389902917e-12 pb0=2.778258873e-17 b1=6.680143798e-10 lb1=-1.335285260e-14 wb1=-8.721742706e-16 pb1=1.743377811e-20 keta=-6.067220295e-01 lketa=1.209030459e-05 wketa=7.417874372e-07 pketa=-1.482749265e-11 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.097533665e-01 lpclm=-7.371783048e-06 wpclm=-6.133801217e-07 ppclm=1.226077551e-11 pdiblc1=0.39 pdiblc2=-1.002496346e-02 lpdiblc2=2.067700979e-07 wpdiblc2=1.345297292e-08 ppdiblc2=-2.689097267e-13 pdiblcb=2.362311511e+00 lpdiblcb=-5.032060181e-05 wpdiblcb=-3.036179439e-06 ppdiblcb=6.068979610e-11 drout=0.56 pscbe1=6.864776709e+08 lpscbe1=2.268208620e+03 wpscbe1=1.323383224e+02 ppscbe1=-2.645293522e-3 pscbe2=3.058498191e-09 lpscbe2=4.731294787e-14 wpscbe2=9.511793143e-15 ppscbe2=-1.901299966e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.140618095e-09 lalpha0=-2.080077982e-14 walpha0=-1.358653878e-15 palpha0=2.715795575e-20 alpha1=1.140618095e-09 lalpha1=-2.080077982e-14 walpha1=-1.358653878e-15 palpha1=2.715795575e-20 beta0=-2.787860768e+02 lbeta0=5.698120552e-03 wbeta0=3.668365471e-04 pbeta0=-7.332648052e-9 agidl=-4.072098903e-08 lagidl=2.755047698e-12 wagidl=2.189357372e-14 pagidl=-4.376277990e-19 bgidl=1000000000.0 cgidl=300.0 egidl=-9.625313682e-02 legidl=1.962312938e-05 pegidl=7.105427358e-27 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.391529389e-01 lkt1=3.965420793e-06 wkt1=2.349112556e-07 pkt1=-4.695610549e-12 kt2=1.798475998e-01 lkt2=-4.641536982e-06 wkt2=-2.796789008e-07 pkt2=5.590465191e-12 at=-7.387347856e+05 lat=1.476647359e+01 wat=9.645083882e-01 pat=-1.927943279e-5 ute=-2.946327405e+00 lute=5.624990520e-05 wute=3.351934983e-06 pute=-6.700139263e-11 ua1=6.923187214e-09 lua1=-1.019524901e-13 wua1=-5.555535708e-15 pua1=1.110488811e-19 ub1=-6.624446708e-18 lub1=1.181053943e-22 wub1=6.139756876e-24 pub1=-1.227268020e-28 uc1=5.276253915e-09 luc1=-1.056414815e-13 wuc1=-6.190964541e-15 puc1=1.237503854e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.061742+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.44751769 k2=0.02149811 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.69603492+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='8.3910929+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0095692 ua=-6.5690804e-10 ub=1.02460111e-18 uc=-7.1776909e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160310.0 a0=1.345571 ags=0.151667 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-0.0018702 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.14095898 pdiblc1=0.39 pdiblc2=0.00031929802 pdiblcb=-0.15511953 drout=0.56 pscbe1=799951250.0 pscbe2=5.4254628e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.2785893 agidl=9.710809773e-8 bgidl=1000000000.0 cgidl=300.0 egidl=0.88544965 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.4407715 kt2=-0.052358472 at=0.0 ute=-0.13226612 ua1=1.8227243e-9 ub1=-7.1588888e-19 uc1=-8.7612717e-12 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-01 pvsat=-1.862645149e-21 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595752e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 ppdiblc2=-6.938893904e-30 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+3 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 wpscbe2=-1.323488980e-29 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 uc1=-1.162365659e-11 luc1=2.286722078e-17 wuc1=-2.584939414e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325658e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 wua=1.654361225e-30 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077653e-03 lketa=-3.715224604e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=2.220446049e-22 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048849e-01 lkt1=2.502969993e-8 kt2=-6.021807946e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-02 wat=-2.328306437e-16 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123885e-18 lub1=2.335179770e-24 wub1=6.162975822e-39 uc1=1.777277470e-11 luc1=-9.439132211e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-08 pk2=-1.110223025e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=-1.058181320e-22 peta0=-3.191891196e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=-6.817463261e-22 petab=7.580741590e-28 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 wute=6.661338148e-22 pute=-8.881784197e-28 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 wub1=6.162975822e-39 pub1=6.162975822e-45 uc1=-1.252175596e-10 luc1=1.899978642e-16 wuc1=1.033975766e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.68 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059394261e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.574548827e-8 k1=5.163379589e-01 lk1=-1.485963682e-10 k2=-3.690874683e-03 lk2=-1.907482336e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.279561642e+00 ldsub=-4.971871951e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.292211523e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.589260317e-8 nfactor='6.870411735e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.183217798e-6 eta0=-4.398980000e-02 leta0=2.610515935e-7 etab=-1.632772774e+00 letab=7.979080824e-7 u0=8.009925096e-03 lu0=8.697852353e-10 ua=-7.759682813e-10 lua=1.274097302e-16 ub=6.727035311e-19 lub=1.823100696e-25 uc=-9.895092236e-11 luc=3.384048354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.004043054e+04 lvsat=-2.630819948e-03 wvsat=-1.164153218e-16 a0=1.693335341e+00 la0=-4.775503818e-7 ags=-3.493192284e-01 lags=7.818591912e-07 pags=-8.881784197e-28 a1=0.0 a2=1.009669841e+00 la2=-9.572104471e-9 b0=0.0 b1=0.0 keta=9.793248020e-03 lketa=-2.322682382e-08 pketa=2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.567025060e+00 lpclm=-7.524585059e-7 pdiblc1=6.637643939e-02 lpdiblc1=-2.707173962e-8 pdiblc2=8.111861681e-04 lpdiblc2=-3.769435660e-10 pdiblcb=-3.034907083e-02 lpdiblcb=5.289535676e-9 drout=1.0 pscbe1=7.729094317e+08 lpscbe1=1.324376613e+1 pscbe2=9.028731239e-09 lpscbe2=1.463768495e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.609000049e+00 lbeta0=1.047440030e-6 agidl=1.226892916e-09 lagidl=-1.147148299e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.213729371e-01 lkt1=-5.704969315e-8 kt2=-6.409955753e-02 lkt2=1.536741214e-8 at=8.783879526e+04 lat=-2.578681467e-2 ute=-1.878857286e+00 lute=8.214518228e-7 ua1=-3.360596897e-09 lua1=2.897579860e-15 wua1=-1.654361225e-30 pua1=-3.308722450e-36 ub1=4.154167712e-18 lub1=-3.223006351e-24 wub1=-3.081487911e-39 pub1=-3.081487911e-45 uc1=3.233299061e-10 luc1=-2.535572683e-16 puc1=-1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.69 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.006609654e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.932239947e-11 k1=4.966170030e-01 lk1=9.492387336e-9 k2=-1.761857806e-02 lk2=6.618088114e-09 wk2=-1.387778781e-23 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.644100980e-01 ldsub=2.576142694e-07 pdsub=2.220446049e-28 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.131984112e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.805956571e-8 nfactor='5.759230761e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.399947553e-7 eta0=0.49 etab=-1.216203250e-03 letab=2.890215328e-10 u0=1.119413334e-02 lu0=-6.868786489e-10 ua=-6.998804391e-11 lua=-2.177228284e-16 ub=4.443627388e-19 lub=2.939390328e-25 uc=-5.818012563e-11 luc=1.390886414e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.047293476e+04 lvsat=1.182384171e-2 a0=8.343866772e-01 la0=-5.763614858e-8 ags=9.847587520e-01 lags=1.296684889e-7 a1=0.0 a2=1.171716763e+00 la2=-8.879198318e-8 b0=0.0 b1=0.0 keta=-4.192784488e-02 lketa=2.058066866e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.557003024e-01 lpclm=2.852782422e-07 wpclm=-1.110223025e-22 ppclm=8.326672685e-29 pdiblc1=-3.690848156e-01 lpdiblc1=1.858122041e-07 wpdiblc1=-2.220446049e-22 ppdiblc1=1.249000903e-28 pdiblc2=-8.705633412e-03 lpdiblc2=4.275544022e-09 wpdiblc2=-1.626303259e-24 ppdiblc2=8.673617380e-31 pdiblcb=1.686604462e-01 lpdiblcb=-9.200024691e-08 wpdiblcb=1.110223025e-22 ppdiblcb=1.110223025e-28 drout=1.488187677e+00 ldrout=-2.386603096e-07 wdrout=3.552713679e-21 pscbe1=8.000276611e+08 lpscbe1=-1.352270444e-02 wpscbe1=-1.907348633e-12 pscbe2=9.493699522e-09 lpscbe2=-8.093219498e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.555599215e+00 lbeta0=9.580609553e-8 agidl=-8.222740835e-10 lagidl=8.870614413e-16 pagidl=-8.271806126e-37 bgidl=7.512236789e+08 lbgidl=1.216192801e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.578143445e-01 lkt1=9.652417683e-9 kt2=-1.325100891e-02 lkt2=-9.490917822e-9 at=-2.296195638e+02 lat=1.726719129e-2 ute=4.373883268e-01 lute=-3.108911698e-07 pute=-2.220446049e-28 ua1=4.741250820e-09 lua1=-1.063170433e-15 ub1=-4.602396930e-18 lub1=1.057815405e-24 uc1=-2.829276611e-10 luc1=4.282386859e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.70 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.954474487e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.938216384e-07 wvth0=-6.820117870e-07 pvth0=1.629121556e-13 k1=-3.489492597e+00 lk1=9.616543876e-07 wk1=3.546109364e-06 pk1=-8.470591438e-13 k2=1.907088917e+00 lk2=-4.531367913e-07 wk2=-1.816732860e-06 pk2=4.339629783e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.480511613e+01 ldsub=-3.342043460e-06 wdsub=-1.683114040e-05 pdsub=4.020454508e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.647456119e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.051127044e-07 wvoff=1.543863634e-06 pvoff=-3.687827062e-13 nfactor='1.502722438e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.853840392e-06 wnfactor=-1.406300595e-05 pnfactor=3.359230231e-12 eta0=6.192648726e+00 leta0=-1.362191701e-06 weta0=-6.415747845e-06 peta0=1.532529688e-12 etab=5.997079623e-01 letab=-1.432537339e-07 wetab=-6.990400796e-07 petab=1.669797038e-13 u0=2.792686040e-02 lu0=-4.683825161e-09 wu0=-1.139728315e-08 pu0=2.722469025e-15 ua=3.242098858e-09 lua=-1.008881027e-15 wua=-2.291349287e-15 pua=5.473346041e-22 ub=4.221177318e-18 lub=-6.082286659e-25 wub=-3.848325001e-24 pub=9.192493931e-31 uc=1.720747195e-10 luc=-4.109211072e-17 wuc=-1.727419421e-16 puc=4.126286772e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.135594555e+05 lvsat=-1.776207355e-01 wvsat=-9.187635236e-01 pvsat=2.194650429e-7 a0=5.590577153e+00 la0=-1.193747368e-06 wa0=-6.732004685e-06 pa0=1.608073959e-12 ags=2.197290171e+00 lags=-1.599688912e-7 a1=0.0 a2=-4.779319936e-01 la2=3.052596153e-07 wa2=2.137669664e-06 pa2=-5.106251527e-13 b0=0.0 b1=0.0 keta=-6.672537229e-02 lketa=7.981452239e-09 wketa=8.840165087e-08 pketa=-2.111650234e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-3.339806916e-01 lpclm=2.323160788e-07 wpclm=1.006957741e-06 ppclm=-2.405319957e-13 pdiblc1=7.463804736e-01 lpdiblc1=-8.063898952e-08 wpdiblc1=-3.639711791e-07 ppdiblc1=8.694179555e-14 pdiblc2=5.420951848e-02 lpdiblc2=-1.075299831e-08 wpdiblc2=-5.456616419e-08 ppdiblc2=1.303421964e-14 pdiblcb=1.638952311e+00 lpdiblcb=-4.432088647e-07 wpdiblcb=-2.395690246e-06 ppdiblcb=5.722585289e-13 drout=-2.702161725e+00 ldrout=7.622884521e-07 wdrout=3.718353858e-06 pdrout=-8.882031860e-13 pscbe1=7.999012102e+08 lpscbe1=1.668263473e-2 pscbe2=-4.273794744e-08 lpscbe2=1.239564132e-14 wpscbe2=6.751190807e-14 ppscbe2=-1.612656948e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=2.672541998e+01 lbeta0=-4.244418991e-06 wbeta0=-2.155412933e-05 pbeta0=5.148634872e-12 agidl=1.437897233e-08 lagidl=-2.744060291e-15 wagidl=-5.891772824e-15 pagidl=1.407367775e-21 bgidl=1.888486861e+09 lbgidl=-1.500387762e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=3.021891950e+00 lkt1=-8.454320248e-07 wkt1=-4.264756830e-06 pkt1=1.018722464e-12 kt2=1.509835437e-01 lkt2=-4.872162540e-08 wkt2=-2.658081083e-07 pkt2=6.349358284e-14 at=6.155641632e+05 lat=-1.298274696e-01 wat=-5.748336360e-01 pat=1.373105106e-7 ute=-1.647000087e+00 lute=1.870066905e-07 wute=-8.208162777e-07 pute=1.960683843e-13 ua1=-4.787079780e-09 lua1=1.212861897e-15 wua1=6.187853319e-15 pua1=-1.478092522e-21 ub1=9.994511496e-18 lub1=-2.428948111e-24 wub1=-1.337773188e-23 pub1=3.195538813e-30 uc1=1.189237198e-10 luc1=-5.316637077e-17 wuc1=-4.520521085e-16 puc1=1.079816871e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.71 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.12e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-2.419170667e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.999899358e-07 wvth0=1.687513389e-06 pvth0=-2.611112600e-13 k1=7.999139645e+00 lk1=-1.076928754e-06 wk1=-9.034693050e-06 pk1=1.406061874e-12 k2=-3.794094283e+00 lk2=5.609252328e-07 wk2=4.693225651e-06 pk2=-7.323563243e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-3.515572503e+01 ldsub=5.607737399e-06 wdsub=4.636773827e-05 pdsub=-7.321585318e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='2.299242537e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.977447370e-07 wvoff=-3.433873646e-06 pvoff=5.193042789e-13 nfactor='-6.950990320e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.257178181e-05 wnfactor=9.413840370e-05 pnfactor=-1.641399492e-11 eta0=-1.077748539e+01 leta0=1.654916441e-06 weta0=1.428422239e-05 peta0=-2.160695313e-12 etab=-7.488466977e-01 letab=9.298088860e-08 wetab=9.428994643e-07 petab=-1.213978937e-13 u0=-1.421014232e-02 lu0=2.676662819e-09 wu0=2.352630614e-08 pu0=-3.494709863e-15 ua=-4.463787585e-09 lua=3.218488872e-16 wua=3.210599943e-15 pua=-4.202129878e-22 ub=-5.868961389e-18 lub=1.205995551e-24 wub=1.006658205e-23 pub=-1.574574323e-30 uc=3.546895544e-10 luc=-7.917143810e-17 wuc=-4.845254772e-16 puc=1.033679714e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.847257995e+06 lvsat=2.990644749e-01 wvsat=2.481589201e+00 pvsat=-3.904651579e-7 a0=-1.425669903e+00 la0=-9.811064619e-09 wa0=2.721634213e-06 pa0=1.280954181e-14 ags=1.25 a1=0.0 a2=1.158116137e+01 la2=-1.905433840e-06 wa2=-1.427060330e-05 pa2=2.487776341e-12 b0=0.0 b1=0.0 keta=2.159744099e+00 lketa=-4.050489423e-07 wketa=-2.881863012e-06 pketa=5.288408101e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.614603622e+00 lpclm=4.937325259e-07 wpclm=3.050762012e-06 ppclm=-6.446280479e-13 pdiblc1=-1.033719298e+01 lpdiblc1=1.971346950e-06 wpdiblc1=1.399836863e-05 ppdiblc1=-2.573833947e-12 pdiblc2=-3.167657868e-01 lpdiblc2=5.711768644e-08 wpdiblc2=4.238352535e-07 ppdiblc2=-7.457410800e-14 pdiblcb=-9.803990370e+00 lpdiblcb=1.639073430e-06 wpdiblcb=1.250654056e-05 ppdiblcb=-2.140010330e-12 drout=2.389245913e+01 ldrout=-4.104114793e-06 wdrout=-3.037020488e-05 pdrout=5.358422564e-12 pscbe1=800000000.0 pscbe2=1.033768946e-07 lpscbe2=-1.351486566e-14 wpscbe2=-1.229186268e-13 ppscbe2=1.764530594e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-4.282785357e+01 lbeta0=8.256165896e-06 wbeta0=6.692908699e-05 pbeta0=-1.077943183e-11 agidl=1.161345881e-08 lagidl=-2.506276518e-15 wagidl=-1.516278731e-14 pagidl=3.272249760e-21 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.051036765e+01 lkt1=1.584700140e-06 wkt1=1.289936734e-05 pkt1=-2.069019366e-12 kt2=-2.441216247e+00 lkt2=4.281857850e-07 wkt2=3.117923581e-06 pkt2=-5.590487809e-13 at=-1.404574883e+06 lat=2.325861534e-01 wat=1.872054201e+00 pat=-3.036695988e-7 ute=9.959223438e+00 lute=-1.951416271e-06 wute=-1.336724976e-05 pute=2.547812014e-12 ua1=2.614271089e-08 lua1=-4.413960513e-15 wua1=-3.357033681e-14 pua1=5.762963953e-21 ub1=-4.076849220e-17 lub1=6.761851236e-24 wub1=5.304316841e-23 pub1=-8.828421735e-30 uc1=3.757067888e-10 luc1=-1.062468534e-16 wuc1=-5.589338911e-16 puc1=1.387182292e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.72 pmos lmin=2.0e-05 lmax=0.0001 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.098247561e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=7.297049227e-7 k1=4.276922968e-01 lk1=3.962872071e-07 wk1=8.881784197e-22 k2=1.868581804e-02 lk2=5.621453833e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-2.092832443e-06 lcit=2.417220556e-10 wcit=-1.694065895e-27 pcit=1.761828530e-31 voff='-1.104059252e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=8.155945326e-6 nfactor='1.222262678e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.658803258e-5 eta0=0.08 etab=-0.07 u0=1.124088892e-02 lu0=-3.341517251e-8 ua=-8.365019490e-10 lua=3.589879299e-15 ub=1.509438192e-18 lub=-9.691345396e-24 uc=-1.141297958e-10 luc=8.465863493e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.012865143e+04 lvsat=2.002511953e+0 a0=1.493590774e+00 la0=-2.958748011e-6 ags=1.037010892e-01 lags=9.587843554e-7 a1=0.0 a2=1.012476349e+00 la2=-4.247162113e-06 wa2=-1.776356839e-21 b0=-1.278607675e-07 lb0=2.555792260e-12 b1=-8.023356901e-11 lb1=1.603778381e-15 keta=2.966561342e-02 lketa=-6.303652749e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.647222096e-02 lpclm=3.146871810e-06 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=1.516490733e-03 lpdiblc2=-2.393052950e-8 pdiblcb=-2.424603954e-01 lpdiblcb=1.745845204e-6 drout=0.56 pscbe1=8.000121807e+08 lpscbe1=-1.217936194e+0 pscbe2=1.121877068e-08 lpscbe2=-1.158016781e-13 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-2.498608750e-11 lalpha0=2.498330655e-15 alpha1=-2.498608750e-11 lalpha1=2.498330655e-15 beta0=3.592705243e+01 lbeta0=-5.926392753e-04 pbeta0=9.094947018e-25 agidl=-2.193825010e-08 lagidl=2.379601971e-12 wagidl=-3.308722450e-30 pagidl=1.058791184e-34 bgidl=1000000000.0 cgidl=300.0 egidl=-9.625313682e-02 legidl=1.962312938e-05 pegidl=1.065814104e-26 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.376199758e-01 lkt1=-6.299540746e-8 kt2=-6.009202116e-02 lkt2=1.545849088e-7 at=8.872762352e+04 lat=-1.773564932e+0 ute=-7.066532693e-02 lute=-1.231330245e-6 ua1=2.157031712e-09 lua1=-6.682427407e-15 ub1=-1.357081407e-18 lub1=1.281671407e-23 uc1=-3.504300659e-11 luc1=5.253421821e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.73 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.061742+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.44751769 k2=0.02149811 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.69603492+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='8.3910929+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0095692 ua=-6.5690804e-10 ub=1.02460111e-18 uc=-7.1776909e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160310.0 a0=1.345571 ags=0.151667 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-0.0018702 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.14095898 pdiblc1=0.39 pdiblc2=0.00031929802 pdiblcb=-0.15511953 drout=0.56 pscbe1=799951250.0 pscbe2=5.4254628e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.2785893 agidl=9.710809773e-8 bgidl=1000000000.0 cgidl=300.0 egidl=0.88544965 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.4407715 kt2=-0.052358472 at=0.0 ute=-0.13226612 ua1=1.8227243e-9 ub1=-7.1588888e-19 uc1=-8.7612717e-12 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.74 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-1 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595752e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-07 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 wpdiblc2=8.673617380e-25 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+03 wpscbe1=-1.907348633e-12 ppscbe1=-7.629394531e-18 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 wpscbe2=1.323488980e-29 ppscbe2=-5.293955920e-35 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 pub1=1.232595164e-44 uc1=-1.162365659e-11 luc1=2.286722078e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.75 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325659e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077653e-03 lketa=-3.715224604e-08 wketa=6.938893904e-24 pketa=2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=2.220446049e-22 ppclm=1.332267630e-27 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048848e-01 lkt1=2.502969993e-8 kt2=-6.021807947e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123885e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.76 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=-1.734723476e-22 peta0=-2.255140519e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=7.424616477e-22 petab=-1.058181320e-27 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 wute=4.440892099e-22 pute=1.554312234e-27 ua1=6.024083757e-09 lua1=-6.382649298e-15 pua1=-6.617444900e-36 ub1=-4.182471934e-18 lub1=5.020846495e-24 uc1=-1.252175596e-10 luc1=1.899978642e-16 wuc1=1.033975766e-31 puc1=-2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.77 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059394261e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.574548827e-8 k1=5.163379589e-01 lk1=-1.485963682e-10 k2=-3.690874683e-03 lk2=-1.907482336e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.279561642e+00 ldsub=-4.971871951e-07 pdsub=-8.881784197e-28 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.292211523e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.589260317e-8 nfactor='6.870411735e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.183217798e-6 eta0=-4.398980000e-02 leta0=2.610515935e-7 etab=-1.632772774e+00 letab=7.979080824e-7 u0=8.009925096e-03 lu0=8.697852353e-10 ua=-7.759682813e-10 lua=1.274097302e-16 ub=6.727035311e-19 lub=1.823100696e-25 uc=-9.895092236e-11 luc=3.384048354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.004043054e+04 lvsat=-2.630819948e-3 a0=1.693335341e+00 la0=-4.775503818e-7 ags=-3.493192284e-01 lags=7.818591912e-7 a1=0.0 a2=1.009669841e+00 la2=-9.572104471e-9 b0=0.0 b1=0.0 keta=9.793248020e-03 lketa=-2.322682382e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.567025060e+00 lpclm=-7.524585059e-7 pdiblc1=6.637643939e-02 lpdiblc1=-2.707173962e-8 pdiblc2=8.111861681e-04 lpdiblc2=-3.769435660e-10 pdiblcb=-3.034907083e-02 lpdiblcb=5.289535676e-9 drout=1.0 pscbe1=7.729094317e+08 lpscbe1=1.324376613e+1 pscbe2=9.028731239e-09 lpscbe2=1.463768495e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.609000049e+00 lbeta0=1.047440030e-6 agidl=1.226892916e-09 lagidl=-1.147148299e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.213729371e-01 lkt1=-5.704969315e-8 kt2=-6.409955753e-02 lkt2=1.536741214e-8 at=8.783879526e+04 lat=-2.578681467e-2 ute=-1.878857286e+00 lute=8.214518228e-7 ua1=-3.360596897e-09 lua1=2.897579860e-15 wua1=3.308722450e-30 pua1=1.654361225e-36 ub1=4.154167712e-18 lub1=-3.223006351e-24 uc1=3.233299061e-10 luc1=-2.535572683e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.78 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.006609654e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.932239946e-11 k1=4.966170030e-01 lk1=9.492387336e-9 k2=-1.761857806e-02 lk2=6.618088114e-09 wk2=-1.387778781e-23 pk2=-3.469446952e-30 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.644100980e-01 ldsub=2.576142694e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.131984112e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.805956571e-8 nfactor='5.759230761e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.399947553e-7 eta0=0.49 etab=-1.216203250e-03 letab=2.890215328e-10 u0=1.119413334e-02 lu0=-6.868786489e-10 ua=-6.998804391e-11 lua=-2.177228284e-16 ub=4.443627388e-19 lub=2.939390328e-25 uc=-5.818012563e-11 luc=1.390886414e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.047293476e+04 lvsat=1.182384171e-2 a0=8.343866772e-01 la0=-5.763614858e-08 wa0=-1.776356839e-21 ags=9.847587520e-01 lags=1.296684889e-7 a1=0.0 a2=1.171716763e+00 la2=-8.879198318e-8 b0=0.0 b1=0.0 keta=-4.192784488e-02 lketa=2.058066866e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.557003024e-01 lpclm=2.852782422e-07 wpclm=3.330669074e-22 ppclm=5.551115123e-29 pdiblc1=-3.690848156e-01 lpdiblc1=1.858122041e-07 wpdiblc1=1.387778781e-22 ppdiblc1=9.020562075e-29 pdiblc2=-8.705633412e-03 lpdiblc2=4.275544022e-09 wpdiblc2=2.059984128e-24 ppdiblc2=-8.944667923e-31 pdiblcb=1.686604462e-01 lpdiblcb=-9.200024691e-8 drout=1.488187677e+00 ldrout=-2.386603096e-7 pscbe1=8.000276611e+08 lpscbe1=-1.352270444e-2 pscbe2=9.493699522e-09 lpscbe2=-8.093219498e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.555599215e+00 lbeta0=9.580609553e-8 agidl=-8.222740835e-10 lagidl=8.870614413e-16 pagidl=-8.271806126e-37 bgidl=7.512236789e+08 lbgidl=1.216192801e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.578143445e-01 lkt1=9.652417683e-9 kt2=-1.325100891e-02 lkt2=-9.490917822e-9 at=-2.296195638e+02 lat=1.726719129e-2 ute=4.373883268e-01 lute=-3.108911698e-07 wute=-4.440892099e-22 pute=1.110223025e-28 ua1=4.741250820e-09 lua1=-1.063170433e-15 ub1=-4.602396930e-18 lub1=1.057815405e-24 uc1=-2.829276611e-10 luc1=4.282386859e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.79 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-7.805529006e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.405749910e-8 k1=-4.472461707e-01 lk1=2.349529836e-7 k2=3.484937124e-01 lk2=-8.083515471e-08 wk2=-1.665334537e-22 pk2=-3.469446952e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.654947035e-01 ldsub=1.071489094e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.229584401e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.127005618e-8 nfactor='2.962416109e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.808036061e-8 eta0=6.885077223e-01 leta0=-4.741753964e-8 etab=-6.25e-6 u0=1.814900519e-02 lu0=-2.348188887e-9 ua=1.276324974e-09 lua=-5.393166190e-16 ub=9.196567555e-19 lub=1.804055510e-25 uc=2.387749767e-11 luc=-5.692240336e-18 wuc=1.090521315e-32 puc=-1.918509721e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.534207143e+04 lvsat=1.066075104e-2 a0=-1.848840900e-01 la0=1.858370596e-7 ags=2.197290171e+00 lags=-1.599688912e-7 a1=0.0 a2=1.355998444e+00 la2=-1.328113483e-7 b0=0.0 b1=0.0 keta=9.115381286e-03 lketa=-1.013462857e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.298994868e-01 lpclm=2.596102059e-8 pdiblc1=4.341255753e-01 lpdiblc1=-6.050661960e-9 pdiblc2=7.396602975e-03 lpdiblc2=4.292028164e-10 pdiblcb=-4.163368351e-01 lpdiblcb=4.773805368e-08 wpdiblcb=8.881784197e-22 drout=4.878551563e-01 ldrout=2.891195681e-10 pscbe1=7.999012102e+08 lpscbe1=1.668263473e-2 pscbe2=1.518126485e-08 lpscbe2=-1.439520925e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.233894147e+00 lbeta0=1.726517851e-7 agidl=9.324355294e-09 lagidl=-1.536663918e-15 bgidl=1.888486861e+09 lbgidl=-1.500387762e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.368900827e-01 lkt1=2.854123928e-8 kt2=-7.705617102e-02 lkt2=5.750221250e-9 at=1.224080320e+05 lat=-1.202726455e-2 ute=-2.351187446e+00 lute=3.552159249e-7 ua1=5.215479907e-10 lua1=-5.521001849e-17 ub1=-1.482392574e-18 lub1=3.125399646e-25 wub1=-7.703719778e-40 uc1=-2.688967816e-10 luc1=3.947231239e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.80 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.0e-06 wmax=1.12e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-9.714350746e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.402015211e-08 wvth0=9.322390042e-13 pvth0=-1.732752644e-19 k1=2.481761779e-01 lk1=1.293473497e-07 wk1=4.892214349e-13 pk1=-9.093158759e-20 k2=2.322757765e-01 lk2=-6.737133359e-08 wk2=1.290675229e-13 pk2=-2.398978061e-20 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=4.623670784e+00 ldsub=-6.735316886e-07 wdsub=-6.354215856e-13 pdsub=1.181058096e-19 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.467146457e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.777196275e-08 wvoff=-1.142791696e-12 pvoff=2.124106926e-19 nfactor='1.125237513e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.509947496e-06 wnfactor=1.153157930e-10 pnfactor=-2.143374646e-17 eta0=1.477115255e+00 leta0=-1.987695053e-07 weta0=-9.719470487e-12 peta0=1.806557979e-18 etab=6.007622203e-02 letab=-1.116752908e-08 wetab=1.112744818e-12 petab=-2.068258792e-19 u0=5.973321629e-03 lu0=-3.214847722e-10 wu0=1.652537224e-14 pu0=-3.071570942e-21 ua=-1.709377372e-09 lua=-3.865667163e-17 wua=-1.198109707e-21 pua=2.226926513e-28 ub=2.767251528e-18 lub=-1.448456153e-25 wub=2.228047492e-29 pub=-4.141271871e-36 uc=-6.099048795e-11 luc=9.509139135e-18 wuc=3.251912996e-22 puc=-6.044330686e-29 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.817247553e+05 lvsat=-3.591988964e-02 wvsat=6.934688892e-08 pvsat=-1.288950618e-14 a0=9.092405073e-01 la0=1.180180203e-09 wa0=1.127111264e-11 pa0=-2.094961706e-18 ags=1.25 a1=0.0 a2=-6.617445391e-01 la2=2.288565339e-07 wa2=-2.834559893e-12 pa2=5.268596475e-19 b0=0.0 b1=0.0 keta=-3.126349108e-01 lketa=4.864885374e-08 wketa=-3.646202202e-12 pketa=6.777196032e-19 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.002677566e+00 lpclm=-5.930076705e-08 wpclm=1.479182934e-12 ppclm=-2.749357311e-19 pdiblc1=1.672174298e+00 lpdiblc1=-2.367758932e-07 wpdiblc1=-1.408078795e-11 ppdiblc1=2.617196056e-18 pdiblc2=4.684698606e-02 lpdiblc2=-6.860232403e-09 wpdiblc2=2.059856486e-13 ppdiblc2=-3.828655251e-20 pdiblcb=9.254714851e-01 lpdiblcb=-1.968581093e-07 wpdiblcb=4.377828398e-11 ppdiblcb=-8.137069644e-18 drout=-2.162511566e+00 ldrout=4.929418876e-07 wdrout=4.216895527e-11 pdrout=-7.837943716e-18 pscbe1=800000000.0 pscbe2=-2.076171126e-09 lpscbe2=1.623203347e-15 wpscbe2=-2.133815779e-19 ppscbe2=3.966123388e-26 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.459132804e+01 lbeta0=-9.916237430e-07 wbeta0=2.568908610e-11 pbeta0=-4.774830444e-18 agidl=-1.395172510e-09 lagidl=3.010800586e-16 wagidl=3.595391044e-19 pagidl=-6.682753334e-26 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=5.561426805e-01 lkt1=-1.903345380e-07 wkt1=-5.662080156e-13 pkt1=1.052410843e-19 kt2=2.336833725e-01 lkt2=-5.142806780e-08 wkt2=1.735882893e-12 pkt2=-3.226485534e-19 at=2.014816580e+05 lat=-2.793545395e-02 wat=-6.360928495e-07 pat=1.182305780e-13 ute=-1.508684514e+00 lute=2.343791916e-07 wute=-3.958932316e-12 pute=7.358467498e-19 ua1=-2.657626559e-09 lua1=5.301452092e-16 wua1=-2.987467220e-20 pua1=5.552805322e-27 ub1=4.737798971e-18 lub1=-8.121439041e-25 wub1=3.427805721e-29 pub1=-6.371262494e-36 uc1=-1.038108343e-10 luc1=1.276143166e-17 wuc1=2.399638041e-21 puc1=-4.460207227e-28 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.81 pmos lmin=2.0e-05 lmax=0.0001 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.098247561e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=7.297049227e-7 k1=4.276922968e-01 lk1=3.962872071e-7 k2=1.868581804e-02 lk2=5.621453833e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-2.092832443e-06 lcit=2.417220556e-10 wcit=1.694065895e-27 pcit=-5.421010862e-32 voff='-1.104059252e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=8.155945326e-6 nfactor='1.222262678e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.658803258e-5 eta0=0.08 etab=-0.07 u0=1.124088892e-02 lu0=-3.341517251e-8 ua=-8.365019490e-10 lua=3.589879299e-15 ub=1.509438192e-18 lub=-9.691345396e-24 uc=-1.141297958e-10 luc=8.465863493e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.012865143e+04 lvsat=2.002511953e+0 a0=1.493590774e+00 la0=-2.958748011e-6 ags=1.037010892e-01 lags=9.587843554e-7 a1=0.0 a2=1.012476349e+00 la2=-4.247162113e-6 b0=-1.278607675e-07 lb0=2.555792260e-12 b1=-8.023356901e-11 lb1=1.603778381e-15 keta=2.966561342e-02 lketa=-6.303652749e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.647222096e-02 lpclm=3.146871810e-06 ppclm=-2.664535259e-27 pdiblc1=0.39 pdiblc2=1.516490733e-03 lpdiblc2=-2.393052950e-8 pdiblcb=-2.424603954e-01 lpdiblcb=1.745845204e-6 drout=0.56 pscbe1=8.000121807e+08 lpscbe1=-1.217936194e+0 pscbe2=1.121877068e-08 lpscbe2=-1.158016781e-13 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-2.498608750e-11 lalpha0=2.498330655e-15 alpha1=-2.498608750e-11 lalpha1=2.498330655e-15 beta0=3.592705243e+01 lbeta0=-5.926392753e-4 agidl=-2.193825010e-08 lagidl=2.379601971e-12 wagidl=-1.985233470e-29 pagidl=2.752857079e-33 bgidl=1000000000.0 cgidl=300.0 egidl=-9.625313682e-02 legidl=1.962312938e-5 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.376199758e-01 lkt1=-6.299540746e-8 kt2=-6.009202116e-02 lkt2=1.545849088e-7 at=8.872762352e+04 lat=-1.773564932e+0 ute=-7.066532693e-02 lute=-1.231330245e-06 wute=2.220446049e-22 ua1=2.157031712e-09 lua1=-6.682427407e-15 wua1=-6.617444900e-30 ub1=-1.357081407e-18 lub1=1.281671407e-23 uc1=-3.504300659e-11 luc1=5.253421821e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.82 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.061742+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.44751769 k2=0.02149811 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.69603492+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='8.3910929+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0095692 ua=-6.5690804e-10 ub=1.02460111e-18 uc=-7.1776909e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=160310.0 a0=1.345571 ags=0.151667 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-0.0018702 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.14095898 pdiblc1=0.39 pdiblc2=0.00031929802 pdiblcb=-0.15511953 drout=0.56 pscbe1=799951250.0 pscbe2=5.4254628e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.2785893 agidl=9.710809773e-8 bgidl=1000000000.0 cgidl=300.0 egidl=0.88544965 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.4407715 kt2=-0.052358472 at=0.0 ute=-0.13226612 ua1=1.8227243e-9 ub1=-7.1588888e-19 uc1=-8.7612717e-12 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.83 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-1 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595753e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 wpdiblc2=-1.734723476e-24 ppdiblc2=6.938893904e-30 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+3 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 wpscbe2=-2.646977960e-29 ppscbe2=-2.117582368e-34 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 pub1=-1.232595164e-44 uc1=-1.162365659e-11 luc1=2.286722078e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.84 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325659e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077653e-03 lketa=-3.715224604e-08 pketa=-2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=4.440892099e-22 ppclm=-3.108624469e-27 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048849e-01 lkt1=2.502969993e-8 kt2=-6.021807947e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123885e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.85 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-08 pk2=-1.110223025e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-06 pdsub=1.776356839e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=5.898059818e-23 peta0=3.920475056e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=-9.367506770e-23 petab=-1.176142517e-27 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 wute=8.881784197e-22 pute=-2.220446049e-27 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 uc1=-1.252175596e-10 luc1=1.899978642e-16 wuc1=-2.067951531e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.86 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059394261e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.574548827e-8 k1=5.163379589e-01 lk1=-1.485963682e-10 k2=-3.690874683e-03 lk2=-1.907482336e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.279561642e+00 ldsub=-4.971871951e-07 pdsub=1.776356839e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.292211523e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.589260317e-8 nfactor='6.870411735e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.183217798e-6 eta0=-4.398980000e-02 leta0=2.610515935e-07 peta0=-4.440892099e-28 etab=-1.632772774e+00 letab=7.979080824e-7 u0=8.009925096e-03 lu0=8.697852353e-10 ua=-7.759682813e-10 lua=1.274097302e-16 ub=6.727035311e-19 lub=1.823100696e-25 uc=-9.895092236e-11 luc=3.384048354e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.004043054e+04 lvsat=-2.630819948e-3 a0=1.693335341e+00 la0=-4.775503818e-7 ags=-3.493192284e-01 lags=7.818591912e-7 a1=0.0 a2=1.009669841e+00 la2=-9.572104471e-9 b0=0.0 b1=0.0 keta=9.793248020e-03 lketa=-2.322682382e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.567025060e+00 lpclm=-7.524585059e-7 pdiblc1=6.637643939e-02 lpdiblc1=-2.707173962e-8 pdiblc2=8.111861681e-04 lpdiblc2=-3.769435660e-10 pdiblcb=-3.034907083e-02 lpdiblcb=5.289535676e-9 drout=1.0 pscbe1=7.729094317e+08 lpscbe1=1.324376613e+1 pscbe2=9.028731239e-09 lpscbe2=1.463768495e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.609000049e+00 lbeta0=1.047440030e-6 agidl=1.226892916e-09 lagidl=-1.147148299e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.213729371e-01 lkt1=-5.704969315e-8 kt2=-6.409955753e-02 lkt2=1.536741214e-8 at=8.783879526e+04 lat=-2.578681467e-2 ute=-1.878857286e+00 lute=8.214518228e-7 ua1=-3.360596897e-09 lua1=2.897579860e-15 pua1=-1.654361225e-36 ub1=4.154167712e-18 lub1=-3.223006351e-24 uc1=3.233299061e-10 luc1=-2.535572683e-16 wuc1=-4.135903063e-31 puc1=-2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.87 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.006609654e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.932239947e-11 k1=4.966170030e-01 lk1=9.492387336e-9 k2=-1.761857806e-02 lk2=6.618088114e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.644100980e-01 ldsub=2.576142694e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.131984112e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.805956571e-8 nfactor='5.759230761e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.399947553e-7 eta0=0.49 etab=-1.216203250e-03 letab=2.890215328e-10 u0=1.119413334e-02 lu0=-6.868786489e-10 ua=-6.998804391e-11 lua=-2.177228284e-16 ub=4.443627388e-19 lub=2.939390328e-25 uc=-5.818012563e-11 luc=1.390886414e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.047293476e+04 lvsat=1.182384171e-2 a0=8.343866772e-01 la0=-5.763614858e-8 ags=9.847587520e-01 lags=1.296684889e-7 a1=0.0 a2=1.171716763e+00 la2=-8.879198318e-8 b0=0.0 b1=0.0 keta=-4.192784488e-02 lketa=2.058066866e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.557003024e-01 lpclm=2.852782422e-07 wpclm=-4.440892099e-22 ppclm=-8.326672685e-29 pdiblc1=-3.690848156e-01 lpdiblc1=1.858122041e-07 wpdiblc1=-2.775557562e-22 ppdiblc1=-2.775557562e-29 pdiblc2=-8.705633412e-03 lpdiblc2=4.275544022e-09 wpdiblc2=-6.722053469e-24 ppdiblc2=1.463672933e-30 pdiblcb=1.686604462e-01 lpdiblcb=-9.200024691e-08 wpdiblcb=-1.110223025e-22 drout=1.488187677e+00 ldrout=-2.386603096e-7 pscbe1=8.000276611e+08 lpscbe1=-1.352270445e-2 pscbe2=9.493699522e-09 lpscbe2=-8.093219498e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.555599215e+00 lbeta0=9.580609553e-8 agidl=-8.222740835e-10 lagidl=8.870614413e-16 bgidl=7.512236789e+08 lbgidl=1.216192801e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.578143445e-01 lkt1=9.652417683e-9 kt2=-1.325100891e-02 lkt2=-9.490917822e-9 at=-2.296195638e+02 lat=1.726719129e-2 ute=4.373883268e-01 lute=-3.108911698e-07 pute=-2.220446049e-28 ua1=4.741250820e-09 lua1=-1.063170433e-15 ub1=-4.602396930e-18 lub1=1.057815405e-24 uc1=-2.829276611e-10 luc1=4.282386859e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.88 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-7.805529006e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.405749910e-8 k1=-4.472461707e-01 lk1=2.349529836e-7 k2=3.484937124e-01 lk2=-8.083515471e-08 wk2=4.440892099e-22 pk2=-5.551115123e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.654947035e-01 ldsub=1.071489094e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.229584401e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.127005618e-8 nfactor='2.962416109e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.808036061e-8 eta0=6.885077223e-01 leta0=-4.741753964e-8 etab=-6.25e-6 u0=1.814900519e-02 lu0=-2.348188887e-9 ua=1.276324974e-09 lua=-5.393166190e-16 ub=9.196567555e-19 lub=1.804055510e-25 uc=2.387749767e-11 luc=-5.692240336e-18 wuc=1.494418099e-32 puc=4.543838814e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.534207143e+04 lvsat=1.066075104e-2 a0=-1.848840900e-01 la0=1.858370596e-7 ags=2.197290171e+00 lags=-1.599688912e-7 a1=0.0 a2=1.355998444e+00 la2=-1.328113483e-7 b0=0.0 b1=0.0 keta=9.115381286e-03 lketa=-1.013462857e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.298994868e-01 lpclm=2.596102059e-8 pdiblc1=4.341255753e-01 lpdiblc1=-6.050661960e-9 pdiblc2=7.396602975e-03 lpdiblc2=4.292028164e-10 pdiblcb=-4.163368351e-01 lpdiblcb=4.773805368e-8 drout=4.878551563e-01 ldrout=2.891195681e-10 pscbe1=7.999012102e+08 lpscbe1=1.668263473e-2 pscbe2=1.518126485e-08 lpscbe2=-1.439520925e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.233894147e+00 lbeta0=1.726517851e-7 agidl=9.324355294e-09 lagidl=-1.536663918e-15 bgidl=1.888486861e+09 lbgidl=-1.500387762e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.368900827e-01 lkt1=2.854123928e-8 kt2=-7.705617102e-02 lkt2=5.750221250e-9 at=1.224080320e+05 lat=-1.202726455e-2 ute=-2.351187446e+00 lute=3.552159249e-7 ua1=5.215479907e-10 lua1=-5.521001849e-17 ub1=-1.482392574e-18 lub1=3.125399646e-25 wub1=-1.540743956e-39 uc1=-2.688967816e-10 luc1=3.947231239e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.89 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=9.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='2.148878608e-03+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.049802015e-07 wvth0=-1.017999868e-06 pvth0=1.892156355e-13 k1=1.181107242e+00 lk1=-4.405654723e-08 wk1=-9.754927563e-07 pk1=1.813148386e-13 k2=-1.189255777e+00 lk2=1.968487362e-07 wk2=1.486384795e-06 pk2=-2.762743418e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=4.828906208e+00 ldsub=-7.116787968e-07 wdsub=-2.145993095e-07 pdsub=3.988757366e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-2.933428059e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.728033849e-07 wvoff=2.391036710e-06 pvoff=-4.444219933e-13 nfactor='-4.835010184e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.568364898e-06 wnfactor=6.232177649e-05 pnfactor=-1.158374860e-11 eta0=1.982978792e+00 leta0=-2.927943610e-07 weta0=-5.289517632e-07 peta0=9.831626422e-14 etab=-3.906706378e-01 letab=7.261278975e-08 wetab=4.713119458e-07 petab=-8.760275136e-14 u0=3.273680204e-03 lu0=1.802975794e-10 wu0=2.822820991e-09 pu0=-5.246777376e-16 ua=2.563693257e-09 lua=-8.328923095e-16 wua=-4.468017855e-15 pua=8.304704788e-22 ub=2.868112101e-18 lub=-1.635925700e-25 wub=-1.054397535e-25 pub=1.959808699e-32 uc=-5.900652882e-11 luc=9.140380651e-18 wuc=-2.074146127e-18 puc=3.855215405e-25 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.188666934e+06 lvsat=-2.044932323e-01 wvsat=-9.483186250e-01 pvsat=1.762639828e-7 a0=7.135228311e+00 la0=-1.156044173e-06 wa0=-6.510018548e-06 pa0=1.210017148e-12 ags=1.250000027e+00 lags=-5.081997045e-15 wags=-2.858905646e-14 pags=5.313847140e-21 a1=0.0 a2=-5.264002574e+00 la2=1.084278235e-06 wa2=4.812219417e-06 pa2=-8.944472230e-13 b0=0.0 b1=0.0 keta=-2.753488950e-01 lketa=4.171850199e-08 wketa=-3.899072461e-08 pketa=7.247205984e-15 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.983923887e-01 lpclm=-5.850428111e-08 wpclm=4.482155003e-09 ppclm=-8.330981505e-16 pdiblc1=2.089114339e+00 lpdiblc1=-3.142725385e-07 wpdiblc1=-4.359757601e-07 ppdiblc1=8.103481453e-14 pdiblc2=7.608195777e-02 lpdiblc2=-1.229413660e-08 wpdiblc2=-3.056852360e-08 ppdiblc2=5.681771482e-15 pdiblcb=-2.781768759e-01 lpdiblcb=2.686401152e-08 wpdiblcb=1.258604985e-06 ppdiblcb=-2.339369085e-13 drout=-2.162471648e+00 ldrout=4.929344682e-07 wdrout=4.305617551e-13 pdrout=-8.002851359e-20 pscbe1=7.999999958e+08 lpscbe1=7.849140167e-07 wpscbe1=4.415588379e-06 ppscbe1=-8.207244873e-13 pscbe2=-2.945237074e-08 lpscbe2=6.711617569e-15 wpscbe2=2.862494321e-14 ppscbe2=-5.320518195e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.807219121e+01 lbeta0=-1.638611781e-06 wbeta0=-3.639641424e-06 pbeta0=6.765001515e-13 agidl=-4.717379679e-08 lagidl=8.809952954e-15 wagidl=4.786749622e-14 pagidl=-8.897131522e-21 bgidl=9.999999970e+08 lbgidl=5.590915680e-07 wbgidl=3.145202637e-06 pbgidl=-5.845985413e-13 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-8.779954171e-01 lkt1=7.622871018e-08 wkt1=1.499565780e-06 pkt1=-2.787242915e-13 kt2=2.336850272e-01 lkt2=-5.142837536e-08 wkt2=5.668548297e-15 pkt2=-1.053613197e-21 at=7.435873295e+05 lat=-1.286966351e-01 wat=-5.668382525e-01 pat=1.053582260e-7 ute=-2.792624130e+00 lute=4.730250480e-07 wute=1.342511550e-06 pute=-2.495326218e-13 ua1=-2.657655258e-09 lua1=5.301505435e-16 wua1=1.340311451e-22 pua1=-2.491237098e-29 ub1=4.737832458e-18 lub1=-8.121501283e-25 wub1=-7.363307315e-31 pub1=1.368617919e-37 uc1=-1.038085303e-10 luc1=1.276100342e-17 wuc1=-9.410079440e-24 puc1=1.749051382e-30 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.90 pmos lmin=2.0e-05 lmax=0.0001 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.180861360e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=8.990165316e-06 wvth0=8.142597765e-08 pvth0=-8.141691494e-12 k1=3.828265016e-01 lk1=4.882367371e-06 wk1=4.422071480e-08 pk1=-4.421579303e-12 k2=1.232146936e-02 lk2=6.925785712e-07 wk2=6.272842076e-09 pk2=-6.272143908e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-2.945947978e-05 lcit=2.978082199e-09 wcit=2.697316969e-11 pcit=-2.697016757e-15 voff='-2.027437464e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.004834893e-04 wvoff=9.101018798e-07 pvoff=-9.100005855e-11 nfactor='2.089356776e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-9.435856231e-04 wnfactor=-8.546270192e-06 pnfactor=8.545318992e-10 eta0=0.08 etab=-0.07 u0=1.502399940e-02 lu0=-4.116841145e-07 wu0=-3.728716917e-09 pu0=3.728301911e-13 ua=-1.242931393e-09 lua=4.422830018e-14 wua=4.005858019e-16 pua=-4.005412167e-20 ub=2.606647261e-18 lub=-1.194000404e-22 wub=-1.081433397e-24 pub=1.081313034e-28 uc=-2.099763664e-10 luc=1.043017664e-14 wuc=9.446848859e-17 puc=-9.445797425e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.665864420e+05 lvsat=2.467149795e+01 wvsat=2.234553838e-01 pvsat=-2.234305132e-5 a0=1.828566468e+00 la0=-3.645258915e-05 wa0=-3.301594137e-07 pa0=3.301226669e-11 ags=-4.848018005e-03 lags=1.181248692e-05 wags=1.069883881e-07 pags=-1.069764803e-11 a1=0.0 a2=1.493320298e+00 la2=-5.232620520e-05 wa2=-4.739303745e-07 pa2=4.738776261e-11 b0=-4.172156850e-07 lb0=3.148806348e-11 wb0=2.851945724e-13 pb0=-2.851628303e-17 b1=-2.618059011e-10 lb1=1.975899069e-14 wb1=1.789616851e-16 pb1=-1.789417666e-20 keta=1.010326392e-01 lketa=-7.766273537e-06 wketa=-7.034091067e-08 pketa=7.033308173e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-3.727464170e-01 lpclm=3.877032609e-05 wpclm=3.511516857e-07 ppclm=-3.511126025e-11 pdiblc1=0.39 pdiblc2=4.225794026e-03 lpdiblc2=-2.948307043e-07 wpdiblc2=-2.670348931e-09 ppdiblc2=2.670051721e-13 pdiblcb=-4.401168727e-01 lpdiblcb=2.150929302e-05 wpdiblcb=1.948145725e-07 ppdiblcb=-1.947928896e-11 drout=0.56 pscbe1=8.001500698e+08 lpscbe1=-1.500530885e+01 wpscbe1=-1.359065045e-01 ppscbe1=1.358913781e-5 pscbe2=2.432929831e-08 lpscbe2=-1.426708520e-12 wpscbe2=-1.292202446e-14 ppscbe2=1.292058623e-18 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-3.078354692e-10 lalpha0=3.078012071e-14 walpha0=2.787825733e-16 palpha0=-2.787515448e-20 alpha1=-3.078354692e-10 lalpha1=3.078012071e-14 walpha1=2.787825733e-16 palpha1=-2.787515448e-20 beta0=1.030229159e+02 lbeta0=-7.301478847e-03 wbeta0=-6.613115916e-05 pbeta0=6.612379877e-9 agidl=-2.913457221e-07 lagidl=2.931735067e-11 wagidl=2.655339314e-13 pagidl=-2.655043775e-17 bgidl=1000000000.0 cgidl=300.0 egidl=-2.317892615e+00 legidl=2.417623504e-04 wegidl=2.189696746e-06 pegidl=-2.189453033e-10 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.304879286e-01 lkt1=-7.761207437e-07 wkt1=-7.029502585e-09 pkt1=7.028720201e-13 kt2=-7.759340585e-02 lkt2=1.904528587e-06 wkt2=1.724974978e-08 pkt2=-1.724782988e-12 at=2.895223996e+05 lat=-2.185080769e+01 wat=-1.979077488e-01 pat=1.978857216e-5 ute=6.874015874e-02 lute=-1.517032723e-05 wute=-1.374011136e-07 pute=1.373858209e-11 ua1=2.913585076e-09 lua1=-8.232934333e-14 wua1=-7.456756393e-16 pua1=7.455926456e-20 ub1=-2.808130188e-18 lub1=1.579054420e-22 wub1=1.430185601e-24 pub1=-1.430026422e-28 uc1=-9.451980607e-11 luc1=6.472360153e-15 wuc1=5.862164205e-17 puc1=-5.861511747e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.91 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-5.109833410e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.399939328e-06 wvth0=-5.428398510e-07 pvth0=4.336677001e-12 k1=7.466229913e-01 lk1=-2.389513369e-06 wk1=-2.948047653e-07 pk1=2.355156945e-12 k2=6.392710121e-02 lk2=-3.389596950e-07 wk2=-4.181894717e-08 pk2=3.340861325e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.924443156e-04 lcit=-1.457523920e-09 wcit=-1.798211312e-10 pcit=1.436567641e-15 voff='5.459819825e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.917832330e-05 wvoff=-6.067345865e-06 pvoff=4.847123736e-11 nfactor='-4.941518031e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.618068019e-04 wnfactor=5.697513461e-05 pnfactor=-4.551669437e-10 eta0=0.08 etab=-0.07 u0=-1.565153653e-02 lu0=2.014851855e-07 wu0=2.485811278e-08 pu0=-1.985882315e-13 ua=2.052621590e-09 lua=-2.164607997e-14 wua=-2.670572013e-15 pua=2.133485263e-20 ub=-6.290126019e-18 lub=5.843640412e-23 wub=7.209555982e-24 pub=-5.759620550e-29 uc=5.672002282e-10 luc=-5.104705282e-15 wuc=-6.297899239e-16 puc=5.031309830e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.671743956e+06 lvsat=-1.207464939e+01 wvsat=-1.489702558e+00 pvsat=1.190104008e-5 a0=-8.876002948e-01 la0=1.784051516e-05 wa0=2.201062758e-06 pa0=-1.758400424e-11 ags=8.753277147e-01 lags=-5.781231374e-06 wags=-7.132559209e-07 pags=5.698108829e-12 a1=0.0 a2=-2.405626326e+00 la2=2.560933198e-05 wa2=3.159535830e-06 pa2=-2.524112101e-11 b0=1.929032783e-06 lb0=-1.541079213e-11 wb0=-1.901297150e-12 pb0=1.518921576e-17 b1=1.210482214e-09 lb1=-9.670385043e-15 wb1=-1.193077901e-15 pb1=9.531344247e-21 keta=-4.776503718e-01 lketa=3.800945941e-06 wketa=4.689394045e-07 pketa=-3.746295940e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.516120287e+00 lpclm=-1.897485491e-05 wpclm=-2.341011238e-06 ppclm=1.870203445e-11 pdiblc1=0.39 pdiblc2=-1.774272394e-02 lpdiblc2=1.442951454e-07 wpdiblc2=1.780232621e-08 ppdiblc2=-1.422204698e-13 pdiblcb=1.162590319e+00 lpdiblcb=-1.052701268e-05 wpdiblcb=-1.298763817e-06 ppdiblcb=1.037565529e-11 drout=0.56 pscbe1=7.990319895e+08 lpscbe1=7.343852554e+00 wpscbe1=9.060433631e-01 ppscbe1=-7.238262642e-6 pscbe2=-8.197805468e-08 lpscbe2=6.982553387e-13 wpscbe2=8.614682971e-14 ppscbe2=-6.882158234e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.985662544e-09 lalpha0=-1.506431293e-14 walpha0=-1.858550488e-15 palpha0=1.484771824e-20 alpha1=1.985662544e-09 lalpha1=-1.506431293e-14 walpha1=-1.858550488e-15 palpha1=1.484771824e-20 beta0=-4.410271673e+02 lbeta0=3.573467540e-03 wbeta0=4.408743944e-04 pbeta0=-3.522088223e-9 agidl=1.893157911e-06 lagidl=-1.434840847e-11 wagidl=-1.770226209e-12 pagidl=1.414210706e-17 bgidl=1000000000.0 cgidl=300.0 egidl=1.569637951e+01 legidl=-1.183225932e-04 wegidl=-1.459797831e-05 pegidl=1.166213510e-10 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.883184811e-01 lkt1=3.798466506e-07 wkt1=4.686335057e-08 pkt1=-3.743852154e-13 kt2=6.431742593e-02 lkt2=-9.321085807e-07 wkt2=-1.149983319e-07 pkt2=9.187067235e-13 at=-1.338631840e+06 lat=1.069415575e+01 wat=1.319384992e+00 pat=-1.054039518e-5 ute=-1.061636024e+00 lute=7.424615349e-06 wute=9.160074240e-07 pute=-7.317864229e-12 ua1=-3.220964791e-09 lua1=4.029337646e-14 wua1=4.971170929e-15 pua1=-3.971403830e-20 ub1=8.957769659e-18 lub1=-7.728160049e-23 wub1=-9.534570676e-24 pub1=7.617044564e-29 uc1=3.877507248e-10 luc1=-3.167682794e-15 wuc1=-3.908109470e-16 puc1=3.122137850e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.92 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 wua=-1.654361225e-30 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-1 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595752e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 wpdiblc2=8.673617380e-25 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+3 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 pub1=1.232595164e-44 uc1=-1.162365659e-11 luc1=2.286722078e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.93 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325658e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077653e-03 lketa=-3.715224604e-08 pketa=2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=3.330669074e-22 ppclm=2.220446049e-28 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 wagidl=3.308722450e-30 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048848e-01 lkt1=2.502969993e-8 kt2=-6.021807946e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123885e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.94 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=5.377642776e-23 peta0=-2.185751580e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=3.920475056e-22 petab=4.631711681e-28 u0=1.292093949e-02 lu0=-3.986569568e-09 wu0=2.775557562e-23 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-02 wat=2.328306437e-16 ute=9.019606480e-01 lute=-1.928415607e-06 wute=-4.440892099e-22 pute=-6.661338148e-28 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 pub1=6.162975822e-45 uc1=-1.252175596e-10 luc1=1.899978642e-16 puc1=-2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.95 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.096500166e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=6.243840458e-08 wvth0=3.657239633e-08 pvth0=-3.616534556e-14 k1=4.467500259e-01 lk1=6.866482286e-08 wk1=6.858739762e-08 pk1=-6.782401988e-14 k2=3.540557254e-02 lk2=-3.885205200e-08 wk2=-3.853431850e-08 pk2=3.810543154e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.912433260e+00 ldsub=-1.123014953e-06 wdsub=-6.237721905e-07 pdsub=6.168296060e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-2.991371208e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.401751929e-06 wvoff=2.328187063e-06 pvoff=-2.302274341e-12 nfactor='-3.639773682e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.209989255e-06 wnfactor=1.035906997e-05 pnfactor=-1.024377352e-11 eta0=-4.574898055e-01 leta0=6.699493440e-07 weta0=4.075547024e-07 peta0=-4.030186186e-13 etab=-1.633094605e+00 letab=7.982263309e-07 wetab=3.172031693e-10 petab=-3.136726980e-16 u0=-3.130902682e-02 lu0=3.975111721e-08 wu0=3.875362402e-08 pu0=-3.832229619e-14 ua=-8.360635370e-09 lua=7.627659475e-15 wua=7.475614746e-15 pua=-7.392411154e-21 ub=2.781703904e-18 lub=-1.903217129e-24 wub=-2.078677165e-24 pub=2.055541488e-30 uc=-1.149161555e-10 luc=4.962802368e-17 wuc=1.573568506e-17 puc=-1.556054688e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.750242027e+05 lvsat=-4.228845227e-01 wvsat=-4.188733555e-01 pvsat=4.142112950e-7 a0=2.034730903e+00 la0=-8.151462117e-07 wa0=-3.364869772e-07 pa0=3.327418771e-13 ags=-3.493192291e-01 lags=7.818591918e-07 wags=6.444036416e-16 pags=-6.372298245e-22 a1=0.0 a2=5.823493325e-01 la2=4.129923269e-07 wa2=4.211764944e-07 pa2=-4.164888000e-13 b0=9.707705920e-16 lb0=-9.599659153e-22 wb0=-9.568128524e-22 pb0=9.461635254e-28 b1=4.035937759e-19 lb1=-3.991017772e-25 wb1=-3.977909046e-25 pb1=3.933634918e-31 keta=4.804604229e-03 lketa=-1.829370363e-08 wketa=4.916917070e-09 pketa=-4.862191783e-15 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.914299633e+00 lpclm=-1.095867913e-06 wpclm=-3.422814592e-07 ppclm=3.384718665e-13 pdiblc1=1.168996606e-01 lpdiblc1=-7.703263734e-08 wpdiblc1=-4.979679830e-08 ppdiblc1=4.924255993e-14 pdiblc2=1.466407932e-03 lpdiblc2=-1.024872712e-09 wpdiblc2=-6.458009852e-10 ppdiblc2=6.386132203e-16 pdiblcb=-2.066815844e-01 lpdiblcb=1.796594684e-07 wpdiblcb=1.737972047e-07 ppdiblcb=-1.718628418e-13 drout=5.811830963e-01 ldrout=4.141554715e-07 wdrout=4.127951542e-07 pdrout=-4.082007441e-13 pscbe1=2.050336954e+08 lpscbe1=5.747990455e+02 wpscbe1=5.597108190e+02 ppscbe1=-5.534812376e-4 pscbe2=6.811211336e-08 lpscbe2=-5.827940723e-14 wpscbe2=-5.823388125e-14 ppscbe2=5.758573815e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.343431244e+00 lbeta0=1.310053054e-06 wbeta0=2.617504563e-07 pbeta0=-2.588371737e-13 agidl=-9.755501537e-09 lagidl=1.074544557e-14 wagidl=1.082448959e-14 pagidl=-1.070401302e-20 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=9.622061795e-02 lkt1=-5.688824319e-07 wkt1=-5.101515949e-07 pkt1=5.044736077e-13 kt2=-8.716677806e-02 lkt2=3.817789451e-08 wkt2=2.273556004e-08 pkt2=-2.248251325e-14 at=1.263791376e+05 lat=-6.389820300e-02 wat=-3.798620930e-02 pat=3.756342279e-8 ute=-1.913227686e+00 lute=8.554396804e-07 wute=3.387622248e-08 pute=-3.349918012e-14 ua1=-4.133738016e-09 lua1=3.662115918e-15 wua1=7.620248955e-16 pua1=-7.535435584e-22 ub1=5.503375746e-18 lub1=-4.557197700e-24 wub1=-1.329809122e-24 pub1=1.315008346e-30 uc1=4.331615978e-10 luc1=-3.621665333e-16 wuc1=-1.082525317e-16 puc1=1.070476810e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.96 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.278311227e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.513203782e-07 wvth0=2.677950480e-07 pvth0=-1.492031633e-13 k1=1.084757674e+00 lk1=-2.432379762e-07 wk1=-5.796843847e-07 pk1=2.490966063e-13 k2=-3.452969821e-01 lk2=1.472620059e-07 wk2=3.229670439e-07 pk2=-1.386217395e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.848905686e+00 ldsub=7.157908182e-07 wdsub=1.561713711e-06 pdsub=-4.515888864e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='3.536360621e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.894603305e-07 wvoff=-4.089896673e-06 pvoff=8.353342551e-13 nfactor='4.123717397e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.272900414e-05 wnfactor=-3.496784134e-05 pnfactor=1.191519361e-11 eta0=1.317000017e+00 leta0=-1.975454955e-07 weta0=-8.151094106e-07 peta0=1.947051863e-13 etab=-1.281599537e-03 letab=4.819070393e-10 wetab=6.445601891e-11 petab=-1.901121986e-16 u0=8.594045236e-02 lu0=-1.756863567e-08 wu0=-7.367161644e-08 pu0=1.663903112e-14 ua=1.420332019e-08 lua=-3.403181479e-15 wua=-1.406808661e-14 pua=3.139658126e-21 ub=-3.440248070e-18 lub=1.138508533e-24 wub=3.828757875e-24 pub=-8.324262797e-31 uc=-3.747081394e-11 luc=1.176731953e-17 wuc=-2.041155320e-17 puc=2.110753484e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-7.477744267e+05 lvsat=1.749050433e-01 wvsat=7.572015009e-01 pvsat=-1.607364200e-7 a0=3.949277881e-01 la0=-1.349566276e-08 wa0=4.331403492e-07 pa0=-4.350583392e-14 ags=7.469353827e-01 lags=2.459331998e-07 wags=2.344039449e-07 pags=-1.145930569e-13 a1=0.0 a2=1.983329918e+00 la2=-2.719050519e-07 wa2=-7.999437809e-07 pa2=1.804802690e-13 b0=-1.941541184e-15 lb0=4.637759426e-22 wb0=1.913625705e-21 pb0=-4.571077721e-28 b1=-8.071875518e-19 lb1=1.928128905e-25 wb1=7.955818092e-25 pb1=-1.900406268e-31 keta=-1.416863263e-02 lketa=-9.018257333e-09 wketa=-2.736009030e-08 pketa=1.091706881e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.265185887e+00 lpclm=4.584871736e-07 wpclm=6.992846010e-07 ppclm=-1.707185333e-13 pdiblc1=-5.151856770e-01 lpdiblc1=2.319749217e-07 wpdiblc1=1.440002233e-07 ppdiblc1=-4.549899001e-14 pdiblc2=-1.668860894e-02 lpdiblc2=7.850570385e-09 wpdiblc2=7.868196303e-09 ppdiblc2=-3.523624634e-15 pdiblcb=-2.523915908e-01 lpdiblcb=2.020057192e-07 wpdiblcb=4.149981508e-07 ppdiblcb=-2.897787484e-13 drout=2.754316326e+00 ldrout=-6.482241706e-07 wdrout=-1.247924252e-06 pdrout=4.036751518e-13 pscbe1=1.935803422e+09 lpscbe1=-2.713223510e+02 wpscbe1=-1.119445577e+03 ppscbe1=2.674079500e-4 pscbe2=-1.120279352e-07 lpscbe2=2.978565831e-14 wpscbe2=1.197743967e-13 ppscbe2=-2.943716867e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.581254503e+00 lbeta0=2.160483970e-07 wbeta0=-2.528641655e-08 pbeta0=-1.185134577e-13 agidl=-1.013064283e-08 lagidl=1.092884090e-14 wagidl=9.174533024e-15 pagidl=-9.897398753e-21 bgidl=5.281633166e+08 lbgidl=2.306667994e+02 wbgidl=2.198532004e+02 pbgidl=-1.074796341e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.803401991e+00 lkt1=-1.403472190e-06 wkt1=-2.327266767e-06 pkt1=1.392806702e-12 kt2=3.472639696e-02 lkt2=-2.141202197e-08 wkt2=-4.728758674e-08 pkt2=1.174970251e-14 at=-1.224106452e+05 lat=5.772765811e-02 wat=1.204243068e-01 pat=-3.987872624e-8 ute=8.255450053e-01 lute=-4.834641252e-07 wute=-3.825757618e-07 pute=1.700917015e-13 ua1=6.337484800e-09 lua1=-1.456950780e-15 wua1=-1.573283328e-15 pua1=3.881185728e-22 ub1=-7.250399985e-18 lub1=1.677740641e-24 wub1=2.609930067e-24 pub1=-6.110119511e-31 uc1=-4.402376540e-10 luc1=6.481215895e-17 wuc1=1.550481898e-16 puc1=-2.167214271e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.97 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-2.110089717e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.036261116e-07 wvth0=-5.613550262e-07 pvth0=4.885591495e-14 k1=2.500047514e+00 lk1=-5.813082601e-07 wk1=-2.904917496e-06 pk1=8.045250396e-13 k2=-1.157335456e+00 lk2=3.412336362e-07 wk2=1.484178357e-06 pk2=-4.160002858e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.734633138e+01 ldsub=4.417660893e-06 wdsub=1.745716545e-05 pdsub=-4.248535442e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='4.004146000e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-9.012002238e-07 wvoff=-4.264889332e-06 pvoff=8.771347517e-13 nfactor='-7.112457618e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.411084711e-05 wnfactor=7.302176951e-05 pnfactor=-1.388028473e-11 eta0=-4.452025897e+00 leta0=1.180501725e-06 weta0=5.066623027e-06 peta0=-1.210264241e-12 etab=-7.447189740e-01 letab=1.780667927e-07 wetab=7.340052444e-07 petab=-1.755065483e-13 u0=3.618763517e-02 lu0=-5.684180229e-09 wu0=-1.777927056e-08 pu0=3.288026459e-15 ua=7.440939352e-09 lua=-1.787851569e-15 wua=-6.075979553e-15 pua=1.230583514e-21 ub=-4.271439599e-18 lub=1.337055253e-24 wub=5.116458771e-24 pub=-1.140019393e-30 uc=3.347570743e-10 luc=-7.714675613e-17 wuc=-3.064097501e-16 puc=7.042714277e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.142545620e+06 lvsat=2.692040382e-01 wvsat=1.151095802e+00 pvsat=-2.548259517e-7 a0=4.891591352e+00 la0=-1.087613688e-06 wa0=-5.003485878e-06 pa0=1.255141073e-12 ags=3.046659586e+00 lags=-3.034019207e-07 wags=-8.371571814e-07 pags=1.413707494e-13 a1=0.0 a2=3.576415423e+00 la2=-6.524453865e-07 wa2=-2.188491824e-06 pa2=5.121627400e-13 b0=0.0 b1=0.0 keta=1.356768448e+00 lketa=-3.364939978e-07 wketa=-1.328276511e-06 pketa=3.216669743e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.097820927e+00 lpclm=4.185087055e-07 wpclm=1.604317049e-06 ppclm=-3.869036343e-13 pdiblc1=-5.701544345e+00 lpdiblc1=1.470840417e-06 wpdiblc1=6.047451258e-06 ppdiblc1=-1.455656339e-12 pdiblc2=-1.347910092e-01 lpdiblc2=3.606169074e-08 wpdiblc2=1.401432387e-07 ppdiblc2=-3.512016401e-14 pdiblcb=-4.372307801e+00 lpdiblcb=1.186130104e-06 wpdiblcb=3.899092016e-06 ppdiblcb=-1.122024250e-12 drout=1.289711006e+01 ldrout=-3.071033310e-06 wdrout=-1.223083464e-05 pdrout=3.027162956e-12 pscbe1=7.998144663e+08 lpscbe1=3.133096612e-02 wpscbe1=8.549668424e-02 ppscbe1=-1.443771768e-8 pscbe2=4.686327011e-08 lpscbe2=-8.168683898e-15 wpscbe2=-3.122648139e-14 ppscbe2=6.632411069e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-1.467118439e+01 lbeta0=5.770358476e-06 wbeta0=2.257574932e-05 pbeta0=-5.517222864e-12 agidl=1.211405757e-07 lagidl=-2.042791508e-14 wagidl=-1.102085268e-13 pagidl=1.861963275e-20 bgidl=2.685132204e+09 lbgidl=-2.845683587e+02 wbgidl=-7.851911759e+02 pbgidl=1.325953161e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.851287320e+01 lkt1=3.449476465e-06 wkt1=1.761896223e-05 pkt1=-3.371749019e-12 kt2=-1.537970646e+00 lkt2=3.542581206e-07 wkt2=1.439909446e-06 pkt2=-3.434970528e-13 at=1.238074386e+04 lat=2.553003901e-02 wat=1.084453158e-01 pat=-3.701730465e-8 ute=1.907099889e+00 lute=-7.418151404e-07 wute=-4.197061680e-06 pute=1.081257953e-12 ua1=1.533516198e-08 lua1=-3.606225928e-15 wua1=-1.460062385e-14 pua1=3.499959402e-21 ub1=-2.462906326e-17 lub1=5.828981938e-24 wub1=2.281386785e-23 pub1=-5.437126570e-30 uc1=-1.307216976e-10 luc1=-9.121917570e-18 wuc1=-1.361884026e-16 puc1=4.789554212e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.98 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.6e-07 wmax=9.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='4.355120427e-03+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.540877883e-07 wvth0=-1.020174389e-06 pvth0=1.390549534e-13 k1=-1.049609291e+01 lk1=1.775764550e-06 wk1=1.053381261e-05 pk1=-1.612340871e-12 k2=6.133871344e+00 lk2=-9.796312703e-07 wk2=-5.731450404e-06 pk2=8.832902352e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=5.324281792e+01 ldsub=-8.258022104e-06 wdsub=-4.793241580e-05 pdsub=7.477729557e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.051158936e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=8.770562406e-07 wvoff=5.463940852e-06 pvoff=-8.428625015e-13 nfactor='8.588042546e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.365114550e-05 wnfactor=-6.997878429e-05 pnfactor=1.130191168e-11 eta0=1.518504107e+01 leta0=-2.350599804e-06 weta0=-1.354119479e-05 peta0=2.126534580e-12 etab=1.523527716e+00 letab=-2.256063863e-07 wetab=-1.415364064e-06 petab=2.063286293e-13 u0=1.319824146e-02 lu0=-1.983363233e-09 wu0=-6.959044920e-09 pu0=1.607873960e-15 ua=-5.049960985e-09 lua=3.538505724e-16 wua=3.036167266e-15 pua=-3.392094139e-22 ub=1.314208153e-17 lub=-1.764995698e-24 wub=-1.023169005e-23 pub=1.597976241e-30 uc=-7.544714579e-10 luc=1.175418525e-16 wuc=6.833913882e-16 puc=-1.064573539e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.498853094e+06 lvsat=-3.805221980e-01 wvsat=-2.239666928e+00 pvsat=3.497620040e-7 a0=-8.134220272e+00 la0=1.224004769e-06 wa0=8.539885903e-06 pa0=-1.135811450e-12 ags=1.249999397e+00 lags=9.398935319e-14 wags=5.923722171e-13 pags=-9.233305676e-20 a1=0.0 a2=-1.062188100e+01 la2=1.920910844e-06 wa2=1.009306226e-05 pa2=-1.719050729e-12 b0=0.0 b1=0.0 keta=-3.899529475e+00 lketa=6.066195312e-07 wketa=3.533081387e-06 pketa=-5.495316762e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.315703600e+00 lpclm=-7.314421811e-07 wpclm=-4.250754756e-06 ppclm=6.624293007e-13 pdiblc1=1.826469387e+01 lpdiblc1=-2.835696021e-06 wpdiblc1=-1.637898281e-05 ppdiblc1=2.566205270e-12 pdiblc2=5.027718896e-01 lpdiblc2=-7.881182538e-08 wpdiblc2=-4.511235076e-07 ppdiblc2=7.124306893e-14 pdiblcb=1.696530174e+01 lpdiblcb=-2.660484668e-06 wpdiblcb=-1.573694690e-05 ppdiblcb=2.414773072e-12 drout=-3.796252626e+01 ldrout=6.073088969e-06 wdrout=3.528532186e-05 pdrout=-5.499923119e-12 pscbe1=7.999999963e+08 lpscbe1=5.753192902e-07 wpscbe1=3.940093994e-06 ppscbe1=-6.141414642e-13 pscbe2=-8.034473494e-08 lpscbe2=1.465313350e-14 wpscbe2=7.878557700e-14 ppscbe2=-1.314785101e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.157188191e+01 lbeta0=-1.153744315e-05 wbeta0=-6.622633357e-05 pbeta0=1.043300613e-11 agidl=1.067426891e-09 lagidl=-1.663798296e-16 wagidl=3.198848485e-16 pagidl=-4.986045133e-23 bgidl=9.999969400e+08 lbgidl=4.769605656e-04 wbgidl=3.016208206e-03 pbgidl=-4.701363716e-10 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=1.553610316e+01 lkt1=-2.531950894e-06 wkt1=-1.467853089e-05 pkt1=2.291954906e-12 kt2=3.968742406e+00 lkt2=-6.336117692e-07 wkt2=-3.681354719e-06 pkt2=5.738127599e-13 at=1.445723757e+06 lat=-2.383153394e-01 wat=-1.258879362e+00 pat=2.134008325e-7 ute=-1.667258710e+01 lute=2.636913378e-06 wute=1.502290841e-05 pute=-2.382308566e-12 ua1=-4.116056328e-08 lua1=6.531598814e-15 wua1=3.794931334e-14 pua1=-5.915159472e-21 ub1=6.372135967e-17 lub1=-1.000591249e-23 wub1=-5.813546279e-23 pub1=9.061574586e-30 uc1=-1.030594110e-09 luc1=1.572190720e-16 wuc1=9.134602471e-16 puc1=-1.423810487e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.99 pmos lmin=2.0e-05 lmax=0.0001 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.100 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.110394410e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.886777775e-7 k1=4.210956021e-01 lk1=2.110826255e-7 k2=1.775005695e-02 lk2=2.994270855e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 pcit=8.131516294e-32 voff='-1.239825132e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.344269313e-6 nfactor='1.349753009e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.079466284e-05 wnfactor=-1.136868377e-19 eta0=0.08 etab=-0.07 u0=1.179712614e-02 lu0=-1.779861227e-8 ua=-8.962599665e-10 lua=1.912151425e-15 ub=1.670762721e-18 lub=-5.162101108e-24 uc=-1.282222813e-10 luc=4.509347416e-16 wuc=8.271806126e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.679434283e+04 lvsat=1.066639228e+0 a0=1.542842824e+00 la0=-1.575978955e-6 ags=8.774092800e-02 lags=5.106970788e-7 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=-1.704051167e-07 lb0=1.361344325e-12 b1=-1.069304601e-10 lb1=8.542535445e-16 keta=4.015882949e-02 lketa=-3.357644528e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 ppclm=-5.329070518e-27 pdiblc1=0.39 pdiblc2=1.914844237e-03 lpdiblc2=-1.274661131e-8 pdiblcb=-2.715221659e-01 lpdiblcb=9.299255256e-07 wpdiblcb=1.776356839e-21 drout=0.56 pscbe1=8.000324548e+08 lpscbe1=-6.487344657e-1 pscbe2=1.314643402e-08 lpscbe2=-6.168183535e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.579227219e+01 lbeta0=-3.156696758e-4 agidl=-6.154969226e-08 lagidl=1.267496459e-12 wagidl=-1.588186776e-28 pagidl=1.270549421e-33 bgidl=1000000000.0 cgidl=300.0 egidl=-4.229045954e-01 legidl=1.045227198e-05 wegidl=-1.776356839e-21 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.365713387e-01 lkt1=-3.355454267e-8 kt2=-6.266527973e-02 lkt2=8.233974711e-8 at=1.182508234e+05 lat=-9.446904559e-1 ute=-5.016829954e-02 lute=-6.558688149e-7 ua1=2.268269050e-09 lua1=-3.559399084e-15 ub1=-1.570431596e-18 lub1=6.826830664e-24 uc1=-4.378798232e-11 luc1=2.798238376e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.101 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-01 pvsat=-7.450580597e-21 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595753e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 ppdiblc2=-4.163336342e-29 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-07 wpdiblcb=1.776356839e-21 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+03 wpscbe1=7.629394531e-12 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 ppscbe2=2.117582368e-34 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 pub1=-4.930380658e-44 uc1=-1.162365659e-11 luc1=2.286722078e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.102 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325658e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077654e-03 lketa=-3.715224604e-08 pketa=5.551115123e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=-1.332267630e-21 ppclm=-4.440892099e-27 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048848e-01 lkt1=2.502969993e-8 kt2=-6.021807946e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292611e-09 lua1=-1.003171333e-15 ub1=-2.832123884e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 puc1=2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.103 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=-2.498001805e-22 peta0=9.922618283e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=-7.147060721e-22 petab=7.910339050e-28 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 pute=1.776356839e-27 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 pub1=2.465190329e-44 uc1=-1.252175596e-10 luc1=1.899978642e-16 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.104 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.056116434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.250414331e-8 k1=5.224851534e-01 lk1=-6.227372655e-9 k2=-7.144540537e-03 lk2=3.224478319e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.223655613e+00 ldsub=-4.419034005e-07 pdsub=-3.552713679e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.205557218e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.404503811e-7 nfactor='7.798850790e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.101323326e-6 eta0=-7.462418332e-03 leta0=2.249307616e-7 etab=-1.632744345e+00 letab=7.978799692e-7 u0=1.148324636e-02 lu0=-2.564877967e-9 ua=-1.059609635e-10 lua=-5.351404061e-16 ub=4.864006036e-19 lub=3.665394455e-25 uc=-9.754060033e-11 luc=3.244585840e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.249860650e+04 lvsat=3.449316359e-2 a0=1.663177455e+00 la0=-4.477281531e-7 ags=-3.493192283e-01 lags=7.818591911e-7 a1=0.0 a2=1.047418086e+00 la2=-4.690021102e-8 b0=-8.575503616e-17 lb0=8.480058261e-23 b1=-3.565229431e-20 lb1=3.525548427e-26 keta=1.023393023e-02 lketa=-2.366260124e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.536347840e+00 lpclm=-7.221227228e-7 pdiblc1=6.191336573e-02 lpdiblc1=-2.265833997e-8 pdiblc2=7.533057929e-04 lpdiblc2=-3.197073994e-10 pdiblcb=-1.477237207e-02 lpdiblcb=-1.011379443e-8 drout=1.036997061e+00 ldrout=-3.658528362e-8 pscbe1=8.230739141e+08 lpscbe1=-3.636238561e+1 pscbe2=3.809477986e-09 lpscbe2=5.307539814e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.632459620e+00 lbeta0=1.024241563e-6 agidl=2.197045537e-09 lagidl=-1.074069652e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.670956386e-01 lkt1=-1.183588529e-8 kt2=-6.206186670e-02 lkt2=1.335240081e-08 wkt2=-4.440892099e-22 at=8.443425409e+04 lat=-2.242016604e-2 ute=-1.875821105e+00 lute=8.184494349e-07 pute=-7.105427358e-27 ua1=-3.292299871e-09 lua1=2.830042980e-15 wua1=-6.617444900e-30 pua1=6.617444900e-36 ub1=4.034982618e-18 lub1=-3.105147788e-24 pub1=1.232595164e-44 uc1=3.136276955e-10 luc1=-2.439630433e-16 wuc1=8.271806126e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.105 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.826083314e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.343176261e-8 k1=4.446623754e-01 lk1=3.181784882e-8 k2=1.132757422e-02 lk2=-5.805984424e-09 wk2=-6.938893904e-24 pk2=-1.040834086e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.244403898e-01 ldsub=2.171402925e-07 pdsub=8.881784197e-28 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-9.797583253e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.329269957e-07 wvoff=7.105427358e-21 nfactor='2.625212974e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.279129933e-7 eta0=4.169452362e-01 leta0=1.745059157e-8 etab=-1.210426333e-03 letab=2.719825911e-10 u0=4.591262030e-03 lu0=8.044064145e-10 ua=-1.330850367e-09 lua=6.367127645e-17 ub=7.875179014e-19 lub=2.193322321e-25 uc=-6.000952568e-11 luc=1.409804193e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.833766079e+04 lvsat=-2.582274881e-3 a0=8.732071908e-01 la0=-6.153539006e-8 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=1.100021230e+00 la2=-7.261631000e-8 b0=1.715100723e-16 lb0=-4.096861098e-23 b1=7.130458861e-20 lb1=-1.703252708e-26 keta=-4.438001254e-02 lketa=3.036516966e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.930264200e-01 lpclm=2.699774716e-07 wpclm=1.776356839e-21 pdiblc1=-3.561786926e-01 lpdiblc1=1.817343246e-07 wpdiblc1=-2.220446049e-22 ppdiblc1=-5.551115123e-29 pdiblc2=-8.000440691e-03 lpdiblc2=3.959736644e-09 wpdiblc2=6.071532166e-24 ppdiblc2=-1.170938346e-29 pdiblcb=2.058549522e-01 lpdiblcb=-1.179718745e-07 wpdiblcb=-4.440892099e-22 ppdiblcb=4.440892099e-28 drout=1.376341573e+00 ldrout=-2.024806355e-7 pscbe1=6.996965507e+08 lpscbe1=2.395310605e+1 pscbe2=2.022856548e-08 lpscbe2=-2.719259489e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.553332902e+00 lbeta0=8.518424213e-8 agidl=0.0 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.663972928e-01 lkt1=1.344837144e-7 kt2=-1.748919269e-02 lkt2=-8.437842332e-9 at=1.056349506e+04 lat=1.369303193e-2 ute=4.030997005e-01 lute=-2.956465794e-07 wute=-1.776356839e-21 ua1=4.600244176e-09 lua1=-1.028385029e-15 ub1=-4.368480081e-18 lub1=1.003053022e-24 uc1=-2.690313562e-10 luc1=4.088148730e-17 wuc1=-1.654361225e-30 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.106 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.308647462e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.967875278e-8 k1=-7.076014787e-01 lk1=3.070591157e-7 k2=4.815142591e-01 lk2=-1.181194778e-07 wk2=-4.440892099e-22 pk2=2.775557562e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.930105641e+00 ldsub=-2.736291180e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.052021965e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.734377323e-8 nfactor='9.507044424e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.215950085e-6 eta0=1.142607435e+00 leta0=-1.558883378e-7 etab=6.577949496e-02 letab=-1.572989991e-08 wetab=2.220446049e-22 petab=1.864827737e-29 u0=1.655552535e-02 lu0=-2.053497164e-9 ua=7.317609614e-10 lua=-4.290246915e-16 ub=1.378223032e-18 lub=7.823049762e-26 uc=-3.584695304e-12 luc=6.198427007e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.285098559e+05 lvsat=-1.217820713e-2 a0=-6.333250901e-01 la0=2.983299759e-7 ags=2.122259360e+00 lags=-1.472984367e-7 a1=0.0 a2=1.159853299e+00 la2=-8.690839645e-8 b0=0.0 b1=0.0 keta=-1.099323509e-01 lketa=1.869500404e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.736875497e-01 lpclm=-8.715494325e-9 pdiblc1=9.761327191e-01 lpdiblc1=-1.365149023e-7 pdiblc2=1.995704097e-02 lpdiblc2=-2.718466999e-9 pdiblcb=-6.687792477e-02 lpdiblcb=-5.282417213e-8 drout=-6.083421450e-01 ldrout=2.716007644e-7 pscbe1=7.999088729e+08 lpscbe1=1.538864396e-2 pscbe2=1.238256912e-08 lpscbe2=-8.450863393e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025726182e+01 lbeta0=-3.218332598e-7 agidl=-5.531627378e-10 lagidl=1.321339832e-16 bgidl=1.818113540e+09 lbgidl=-1.381548262e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=9.422220074e-01 lkt1=-2.736541778e-7 kt2=5.199674285e-02 lkt2=-2.503594776e-8 at=1.321275210e+05 lat=-1.534496695e-2 ute=-2.727352100e+00 lute=4.521244422e-7 ua1=-7.870433631e-10 lua1=2.584763459e-16 pua1=-8.271806126e-37 ub1=5.623166473e-19 lub1=-1.747663926e-25 uc1=-2.811027645e-10 luc1=4.376498461e-17 wuc1=1.654361225e-30 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.107 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=8.6e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-9.931543892e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.451509486e-08 wvth0=-1.168078314e-07 pvth0=2.171107163e-14 k1=2.232319638e+00 lk1=-2.084726409e-07 wk1=-9.933178159e-07 pk1=1.846279824e-13 k2=8.272327637e-01 lk2=-1.942691642e-07 wk2=-9.256417598e-07 pk2=1.720490339e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=5.564914671e-01 ldsub=-4.586146319e-08 wdsub=-2.185194647e-07 pdsub=4.061621291e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='1.276215319e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.429054131e-06 wvoff=-1.157380850e-05 pvoff=2.151223786e-12 nfactor='2.876851303e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.304331957e-05 wnfactor=-2.527375647e-04 pnfactor=4.697633115e-11 eta0=8.167465371e-01 leta0=-1.110137198e-07 weta0=-5.289511586e-07 peta0=9.831615184e-14 etab=-5.692749632e-01 letab=1.007241565e-07 wetab=4.799240839e-07 petab=-8.920348947e-14 u0=5.504977956e-02 lu0=-9.415148015e-09 wu0=-4.486071856e-08 pu0=8.338261758e-15 ua=3.236330670e-09 lua=-9.377386158e-16 wua=-4.468080755e-15 pua=8.304821699e-22 ub=1.960605889e-18 lub=-2.214160605e-26 wub=-1.054997168e-25 pub=1.960923236e-32 uc=2.470670693e-12 luc=-4.432691369e-19 wuc=-2.112056181e-18 puc=3.925678823e-25 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.329713827e+06 lvsat=2.576358591e-01 wvsat=1.227567504e+00 pvsat=-2.281679719e-7 a0=8.484088001e+00 la0=-1.366290969e-06 wa0=-6.510019672e-06 pa0=1.210017356e-12 ags=1.249999978e+00 lags=5.733106434e-15 wags=6.674690667e-14 pags=-1.240625380e-20 a1=0.0 a2=-4.887798307e+00 la2=1.028419613e-06 wa2=4.900150830e-06 pa2=-9.107910348e-13 b0=0.0 b1=0.0 keta=4.480033014e-02 lketa=-8.183149155e-09 wketa=-3.899045977e-08 pketa=7.247156758e-15 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.169231343e-01 lpclm=9.579261270e-10 wpclm=4.564207222e-09 ppclm=-8.483491964e-16 pdiblc1=6.690069315e-01 lpdiblc1=-9.317227188e-08 wpdiblc1=-4.439416121e-07 ppdiblc1=8.251542744e-14 pdiblc2=3.900619837e-02 lpdiblc2=-6.532799657e-09 wpdiblc2=-3.112709477e-08 ppdiblc2=5.785593105e-15 pdiblcb=-1.826808881e+00 lpdiblcb=2.689764300e-07 wpdiblcb=1.281601909e-06 ppdiblcb=-2.382113468e-13 drout=1.000002240e+00 ldrout=-3.873937047e-13 wdrout=-1.128322708e-12 pdrout=2.097213425e-19 pscbe1=8.000000120e+08 lpscbe1=-2.218666077e-06 wpscbe1=-1.030905151e-05 ppscbe1=1.916145325e-12 pscbe2=-2.553424115e-08 lpscbe2=6.117437060e-15 wpscbe2=2.914798799e-14 ppscbe2=-5.417736528e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.253625129e+01 lbeta0=-7.778277127e-07 wbeta0=-3.706147693e-06 pbeta0=6.888616717e-13 agidl=5.417498026e-08 lagidl=-1.002688414e-14 wagidl=-4.777548385e-14 pagidl=8.880029183e-21 bgidl=1.000000279e+09 lbgidl=-4.367739868e-05 wbgidl=-7.342895508e-06 pbgidl=1.364822388e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.997128238e-01 lkt1=-5.177728528e-08 wkt1=-2.467053451e-07 pkt1=4.585512250e-14 kt2=-9.625899344e-02 lkt2=-1.726053078e-15 wkt2=-2.076593475e-14 pkt2=3.859764064e-21 at=6.929996725e+05 lat=-1.211390386e-01 wat=-5.771958716e-01 pat=1.072833967e-7 ute=-1.593596795e+00 lute=2.869083286e-07 wute=1.367043055e-06 pute=-2.540922926e-13 ua1=7.435796928e-10 lua1=3.355629547e-23 wua1=-4.230078833e-22 pua1=7.862447675e-29 ub1=-4.726027072e-19 lub1=4.829925600e-31 wub1=1.801473603e-30 pub1=-3.348398998e-37 uc1=-2.193903712e-11 luc1=6.556618174e-24 wuc1=2.276894790e-23 puc1=-4.232064257e-30 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.108 pmos lmin=2.0e-05 lmax=0.0001 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.109 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.110394410e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.886777775e-7 k1=4.210956021e-01 lk1=2.110826255e-7 k2=1.775005695e-02 lk2=2.994270855e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=3.388131789e-27 pcit=3.794707604e-31 voff='-1.239825132e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.344269313e-6 nfactor='1.349753009e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.079466284e-5 eta0=0.08 etab=-0.07 u0=1.179712614e-02 lu0=-1.779861227e-8 ua=-8.962599665e-10 lua=1.912151425e-15 wua=6.617444900e-30 ub=1.670762721e-18 lub=-5.162101108e-24 uc=-1.282222813e-10 luc=4.509347416e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.679434283e+04 lvsat=1.066639228e+0 a0=1.542842824e+00 la0=-1.575978955e-6 ags=8.774092800e-02 lags=5.106970788e-7 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-06 wa2=7.105427358e-21 b0=-1.704051168e-07 lb0=1.361344325e-12 b1=-1.069304601e-10 lb1=8.542535445e-16 keta=4.015882949e-02 lketa=-3.357644528e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 wpclm=1.110223025e-22 ppclm=-6.217248938e-27 pdiblc1=0.39 pdiblc2=1.914844237e-03 lpdiblc2=-1.274661131e-8 pdiblcb=-2.715221659e-01 lpdiblcb=9.299255256e-7 drout=0.56 pscbe1=8.000324548e+08 lpscbe1=-6.487344658e-1 pscbe2=1.314643402e-08 lpscbe2=-6.168183535e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.579227219e+01 lbeta0=-3.156696758e-4 agidl=-6.154969226e-08 lagidl=1.267496459e-12 wagidl=1.191140082e-28 pagidl=-2.329340605e-33 bgidl=1000000000.0 cgidl=300.0 egidl=-4.229045954e-01 legidl=1.045227198e-05 wegidl=8.881784197e-22 pegidl=-2.131628207e-26 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.365713387e-01 lkt1=-3.355454267e-08 wkt1=-3.552713679e-21 kt2=-6.266527973e-02 lkt2=8.233974711e-8 at=1.182508234e+05 lat=-9.446904559e-1 ute=-5.016829954e-02 lute=-6.558688149e-7 ua1=2.268269050e-09 lua1=-3.559399084e-15 ub1=-1.570431596e-18 lub1=6.826830664e-24 uc1=-4.378798232e-11 luc1=2.798238376e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.110 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-1 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595753e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 ppdiblc2=-2.775557562e-29 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+3 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 wpscbe2=-5.293955920e-29 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 uc1=-1.162365659e-11 luc1=2.286722078e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.111 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325658e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077654e-03 lketa=-3.715224604e-08 pketa=5.551115123e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=-1.332267630e-21 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048848e-01 lkt1=2.502969993e-8 kt2=-6.021807946e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123884e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 puc1=-1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.112 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-08 pk2=-2.220446049e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-06 pdsub=3.552713679e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=-2.775557562e-22 peta0=3.469446952e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=-5.412337245e-22 petab=2.116362641e-27 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 wute=-3.552713679e-21 pute=5.329070518e-27 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 uc1=-1.252175596e-10 luc1=1.899978642e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.113 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.056116434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.250414331e-8 k1=5.224851534e-01 lk1=-6.227372655e-9 k2=-7.144540537e-03 lk2=3.224478319e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.223655613e+00 ldsub=-4.419034005e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.205557218e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.404503811e-7 nfactor='7.798850790e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.101323326e-6 eta0=-7.462418332e-03 leta0=2.249307616e-7 etab=-1.632744345e+00 letab=7.978799692e-7 u0=1.148324636e-02 lu0=-2.564877967e-9 ua=-1.059609635e-10 lua=-5.351404061e-16 ub=4.864006036e-19 lub=3.665394455e-25 uc=-9.754060033e-11 luc=3.244585840e-17 wuc=-8.271806126e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.249860650e+04 lvsat=3.449316359e-2 a0=1.663177455e+00 la0=-4.477281531e-7 ags=-3.493192283e-01 lags=7.818591911e-7 a1=0.0 a2=1.047418086e+00 la2=-4.690021102e-8 b0=-8.575503616e-17 lb0=8.480058261e-23 b1=-3.565229431e-20 lb1=3.525548427e-26 keta=1.023393023e-02 lketa=-2.366260124e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.536347840e+00 lpclm=-7.221227228e-7 pdiblc1=6.191336573e-02 lpdiblc1=-2.265833997e-8 pdiblc2=7.533057929e-04 lpdiblc2=-3.197073994e-10 pdiblcb=-1.477237207e-02 lpdiblcb=-1.011379443e-8 drout=1.036997061e+00 ldrout=-3.658528362e-8 pscbe1=8.230739141e+08 lpscbe1=-3.636238561e+1 pscbe2=3.809477986e-09 lpscbe2=5.307539814e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.632459620e+00 lbeta0=1.024241563e-6 agidl=2.197045537e-09 lagidl=-1.074069652e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.670956386e-01 lkt1=-1.183588529e-8 kt2=-6.206186670e-02 lkt2=1.335240081e-8 at=8.443425409e+04 lat=-2.242016604e-2 ute=-1.875821105e+00 lute=8.184494349e-7 ua1=-3.292299871e-09 lua1=2.830042980e-15 wua1=-6.617444900e-30 ub1=4.034982618e-18 lub1=-3.105147788e-24 pub1=6.162975822e-45 uc1=3.136276955e-10 luc1=-2.439630433e-16 wuc1=-8.271806126e-31 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.114 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.826083314e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.343176261e-8 k1=4.446623754e-01 lk1=3.181784882e-8 k2=1.132757422e-02 lk2=-5.805984424e-09 wk2=-2.081668171e-23 pk2=-1.214306433e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.244403898e-01 ldsub=2.171402925e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-9.797583253e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.329269957e-7 nfactor='2.625212974e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.279129933e-7 eta0=4.169452362e-01 leta0=1.745059157e-8 etab=-1.210426333e-03 letab=2.719825911e-10 u0=4.591262030e-03 lu0=8.044064145e-10 ua=-1.330850367e-09 lua=6.367127645e-17 ub=7.875179014e-19 lub=2.193322321e-25 uc=-6.000952568e-11 luc=1.409804193e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.833766079e+04 lvsat=-2.582274881e-3 a0=8.732071908e-01 la0=-6.153539006e-8 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=1.100021230e+00 la2=-7.261631000e-8 b0=1.715100723e-16 lb0=-4.096861098e-23 b1=7.130458861e-20 lb1=-1.703252708e-26 keta=-4.438001254e-02 lketa=3.036516966e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.930264200e-01 lpclm=2.699774716e-07 wpclm=-1.776356839e-21 ppclm=-8.881784197e-28 pdiblc1=-3.561786926e-01 lpdiblc1=1.817343246e-07 wpdiblc1=-6.661338148e-22 ppdiblc1=3.330669074e-28 pdiblc2=-8.000440691e-03 lpdiblc2=3.959736644e-09 wpdiblc2=-2.428612866e-23 ppdiblc2=-1.062518129e-29 pdiblcb=2.058549522e-01 lpdiblcb=-1.179718745e-07 ppdiblcb=-4.440892099e-28 drout=1.376341573e+00 ldrout=-2.024806355e-7 pscbe1=6.996965507e+08 lpscbe1=2.395310605e+1 pscbe2=2.022856548e-08 lpscbe2=-2.719259489e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.553332902e+00 lbeta0=8.518424213e-8 agidl=0.0 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.663972928e-01 lkt1=1.344837144e-7 kt2=-1.748919269e-02 lkt2=-8.437842332e-9 at=1.056349506e+04 lat=1.369303193e-2 ute=4.030997005e-01 lute=-2.956465794e-07 pute=8.881784197e-28 ua1=4.600244176e-09 lua1=-1.028385029e-15 ub1=-4.368480081e-18 lub1=1.003053022e-24 uc1=-2.690313562e-10 luc1=4.088148730e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.115 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='2.168233035e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.660732397e-07 wvth0=-2.656066975e-06 pvth0=6.344547183e-13 k1=-1.023469066e+00 lk1=3.825104063e-07 wk1=2.797392848e-07 pk1=-6.682132296e-14 k2=-1.230143196e+00 lk2=2.907441384e-07 wk2=1.515881498e-06 pk2=-3.620986135e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.935836715e+00 ldsub=-5.138680996e-07 wdsub=-8.906975653e-07 pdsub=2.127609274e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.669242681e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.491974124e-06 wvoff=5.281885462e-06 pvoff=-1.261683980e-12 nfactor='-9.977938716e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.488929983e-05 wnfactor=9.678646811e-05 pnfactor=-2.311938364e-11 eta0=3.379817246e+00 leta0=-6.902906454e-07 weta0=-1.981322228e-06 peta0=4.732784405e-13 etab=2.804513364e-01 letab=-6.700856268e-08 wetab=-1.901181056e-07 petab=4.541351189e-14 u0=9.309045671e-03 lu0=-3.225305638e-10 wu0=6.417641823e-09 pu0=-1.532982102e-15 ua=-1.075622216e-09 lua=2.704928080e-18 wua=1.600658304e-15 pua=-3.823492491e-22 ub=3.218834943e-18 lub=-3.614364695e-25 wub=-1.630086402e-24 pub=3.893787388e-31 uc=-1.122147664e-10 luc=2.656830778e-17 wuc=9.620518080e-17 puc=-2.298053154e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.357470014e+05 lvsat=-6.168094407e-02 wvsat=-1.835337753e-01 pvsat=4.384071290e-8 a0=-2.751867379e+00 la0=8.043861723e-07 wa0=1.876227659e-06 pa0=-4.481745008e-13 ags=2.122259388e+00 lags=-1.472984433e-07 wags=-2.419574230e-14 pags=5.779632772e-21 a1=0.0 a2=1.997655719e+00 la2=-2.870342606e-07 wa2=-7.419762549e-07 pa2=1.772358680e-13 b0=0.0 b1=0.0 keta=-2.201734676e-01 lketa=4.502829959e-08 wketa=9.763195825e-08 pketa=-2.332134587e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.631235178e-01 lpclm=-6.192064035e-09 wpclm=9.355739020e-09 ppclm=-2.234805380e-15 pdiblc1=2.492799844e+00 lpdiblc1=-4.988011784e-07 wpdiblc1=-1.343193772e-06 ppdiblc1=3.208486964e-13 pdiblc2=-1.269330109e-03 lpdiblc2=2.351876259e-09 wpdiblc2=1.879854120e-08 ppdiblc2=-4.490407537e-15 pdiblcb=-6.214551482e+00 lpdiblcb=1.415670610e-06 wpdiblcb=5.444514951e-06 ppdiblcb=-1.300531286e-12 drout=-6.083433780e-01 ldrout=2.716010589e-07 wdrout=1.091991919e-12 pdrout=-2.608441108e-19 pscbe1=7.999088766e+08 lpscbe1=1.538776180e-02 wpscbe1=-3.270675659e-06 ppscbe1=7.812652588e-13 pscbe2=-5.619405608e-09 lpscbe2=3.455045365e-15 wpscbe2=1.594294487e-14 ppscbe2=-3.808291240e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.027741067e+01 lbeta0=-3.266462140e-07 wbeta0=-1.784425886e-08 pbeta0=4.262458114e-15 agidl=-2.449465451e-08 lagidl=5.851038123e-15 wagidl=2.120311183e-14 pagidl=-5.064787322e-21 bgidl=1.818113554e+09 lbgidl=-1.381548295e+02 wbgidl=-1.213946533e-05 pbgidl=2.899753571e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=2.161357738e+01 lkt1=-5.211420835e-06 wkt1=-1.830700708e-05 pkt1=4.372994782e-12 kt2=4.201323668e-01 lkt2=-1.129725043e-07 wkt2=-3.260290076e-07 pkt2=7.787854904e-14 at=-5.390357964e+04 lat=2.909228206e-02 wat=1.647532354e-01 pat=-3.935460534e-8 ute=-6.234815451e+00 lute=1.289952213e-06 wute=3.106286707e-06 pute=-7.419987058e-13 ua1=-3.973509631e-09 lua1=1.019627543e-15 wua1=2.822004629e-15 pua1=-6.740922457e-22 ub1=3.466488140e-18 lub1=-8.684858370e-25 wub1=-2.571998166e-24 pub1=6.143732019e-31 uc1=-3.407032927e-10 luc1=5.800176276e-17 wuc1=5.278353894e-17 puc1=-1.260840395e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.116 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.2e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-6.782500801e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=8.204797135e-07 wvth0=5.010364716e-06 pvth0=-7.266349205e-13 k1=1.241650052e+00 lk1=-2.851902678e-13 wk1=-1.159590357e-07 pk1=2.778285619e-19 k2=2.953107055e+00 lk2=-4.575276194e-07 wk2=-2.808362802e-06 pk2=4.051965135e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.071503902e-01 ldsub=1.246905478e-12 wdsub=3.692163642e-07 pdsub=-8.121330382e-19 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='6.381568141e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.835843113e-07 wvoff=-5.923022010e-06 pvoff=6.939595129e-13 nfactor='2.730174151e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.774315194e-06 wnfactor=-2.213630715e-05 pnfactor=-3.342616188e-12 eta0=-7.078861471e-01 leta0=-1.908779499e-13 weta0=8.212970885e-07 peta0=1.283245954e-19 etab=-1.163551493e-01 letab=1.635138200e-13 wetab=7.880833243e-08 petab=-1.053403134e-19 u0=-2.509519426e-02 lu0=6.039716633e-09 wu0=2.611743345e-08 pu0=-5.348906382e-15 ua=-1.059671604e-09 lua=1.249060394e-20 wua=-6.634466295e-16 pua=-1.084047267e-26 ub=1.078507955e-18 lub=6.041441199e-31 wub=6.757056197e-25 pub=-3.961149418e-37 uc=4.511518326e-11 luc=-9.001619704e-25 wuc=-3.987897469e-17 puc=-2.200399853e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.381677163e+05 lvsat=-6.834025079e-02 wvsat=-2.495450847e-01 pvsat=6.052364245e-8 a0=2.011474541e+00 la0=6.849440410e-13 wa0=-7.777307944e-07 pa0=-5.909088330e-19 ags=1.249999985e+00 lags=2.209453953e-15 wags=5.998725783e-14 pags=-9.285635372e-21 a1=0.0 a2=2.979207143e-01 la2=-1.129221872e-14 wa2=3.075639787e-07 pa2=9.650872101e-21 b0=0.0 b1=0.0 keta=4.647176683e-02 lketa=-8.932938632e-14 wketa=-4.047072088e-08 pketa=5.894958298e-20 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.264555378e-01 lpclm=6.356443194e-14 wpclm=-3.877899051e-09 ppclm=-4.503795026e-20 pdiblc1=-4.609599909e-01 lpdiblc1=2.695344090e-13 wpdiblc1=5.567819536e-07 ppdiblc1=-2.250310684e-19 pdiblc2=1.265778096e-02 lpdiblc2=5.518142804e-15 wpdiblc2=-7.792356648e-09 ppdiblc2=-2.880564148e-21 pdiblcb=2.168643790e+00 lpdiblcb=4.676120611e-13 wpdiblcb=-2.256858877e-06 ppdiblcb=-3.170625238e-19 drout=1.000004036e+00 ldrout=-6.261631498e-13 wdrout=-2.718649313e-12 pdrout=4.211808147e-19 pscbe1=7.999999866e+08 lpscbe1=2.216106415e-06 wpscbe1=1.217721558e-05 ppscbe1=-2.011379242e-12 pscbe2=1.484038863e-08 lpscbe2=-9.757385448e-23 wpscbe2=-6.608672385e-15 ppscbe2=4.017563031e-28 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.343098775e+00 lbeta0=1.139656035e-12 wbeta0=7.400419436e-09 pbeta0=-6.721896284e-19 agidl=1.015352597e-08 lagidl=-1.271299343e-22 wagidl=-8.789115460e-15 pagidl=1.100464676e-28 bgidl=1.000000297e+09 lbgidl=-4.814885712e-05 wbgidl=-2.361618042e-05 pbgidl=5.324844360e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.879941798e+01 lkt1=7.351613286e-06 wkt1=4.261713833e-05 pkt1=-6.510750442e-12 kt2=-2.488580142e-01 lkt2=-1.085374475e-13 wkt2=1.351450292e-07 pkt2=9.845428472e-20 at=1.183725023e+05 lat=2.212370769e-08 wat=-6.829340789e-02 pat=-2.056943020e-14 ute=1.403913598e+00 lute=4.218140015e-14 wute=-1.287618094e-06 pute=-2.156912648e-21 ua1=2.064428120e-09 lua1=1.095570711e-21 wua1=-1.169772848e-15 pua1=-8.619188631e-28 ub1=-1.676437835e-18 lub1=7.956157116e-32 wub1=1.066144675e-24 pub1=2.244745922e-38 uc1=2.766521061e-12 luc1=1.686011016e-23 wuc1=-2.187976307e-17 puc1=-1.335706324e-29 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.117 pmos lmin=2.0e-05 lmax=0.0001 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.118 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.110394410e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.886777775e-7 k1=4.210956021e-01 lk1=2.110826255e-7 k2=1.775005695e-02 lk2=2.994270855e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 pcit=-1.897353802e-31 voff='-1.239825132e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.344269313e-6 nfactor='1.349753009e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.079466284e-5 eta0=0.08 etab=-0.07 u0=1.179712614e-02 lu0=-1.779861227e-8 ua=-8.962599665e-10 lua=1.912151425e-15 ub=1.670762721e-18 lub=-5.162101108e-24 uc=-1.282222813e-10 luc=4.509347416e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.679434283e+04 lvsat=1.066639228e+0 a0=1.542842824e+00 la0=-1.575978955e-6 ags=8.774092800e-02 lags=5.106970788e-7 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=-1.704051167e-07 lb0=1.361344325e-12 b1=-1.069304601e-10 lb1=8.542535445e-16 keta=4.015882949e-02 lketa=-3.357644528e-07 pketa=8.881784197e-28 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=1.914844237e-03 lpdiblc2=-1.274661131e-8 pdiblcb=-2.715221659e-01 lpdiblcb=9.299255256e-7 drout=0.56 pscbe1=8.000324548e+08 lpscbe1=-6.487344658e-1 pscbe2=1.314643402e-08 lpscbe2=-6.168183535e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.579227219e+01 lbeta0=-3.156696758e-4 agidl=-6.154969226e-08 lagidl=1.267496459e-12 wagidl=2.646977960e-29 pagidl=-8.470329473e-34 bgidl=1000000000.0 cgidl=300.0 egidl=-4.229045954e-01 legidl=1.045227198e-05 pegidl=-7.105427358e-27 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.365713387e-01 lkt1=-3.355454267e-8 kt2=-6.266527973e-02 lkt2=8.233974711e-8 at=1.182508234e+05 lat=-9.446904559e-1 ute=-5.016829954e-02 lute=-6.558688149e-7 ua1=2.268269050e-09 lua1=-3.559399084e-15 ub1=-1.570431596e-18 lub1=6.826830664e-24 uc1=-4.378798232e-11 luc1=2.798238376e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.119 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-01 pvsat=-3.725290298e-21 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595752e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-08 wpdiblc2=-1.734723476e-24 ppdiblc2=6.938893904e-30 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+3 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 ppscbe2=2.117582368e-34 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-6 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 uc1=-1.162365659e-11 luc1=2.286722078e-17 wuc1=-5.169878828e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.120 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325658e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077653e-03 lketa=-3.715224604e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=8.881784197e-22 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048849e-01 lkt1=2.502969993e-8 kt2=-6.021807946e-02 lkt2=1.562472077e-8 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123884e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.121 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-06 pdsub=1.776356839e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=-3.434752482e-22 peta0=-1.838806885e-28 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=1.543903894e-21 petab=3.268219029e-27 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767845e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 wute=-8.881784197e-22 pute=-1.332267630e-27 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 pub1=-1.232595164e-44 uc1=-1.252175596e-10 luc1=1.899978642e-16 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.122 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.056116434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.250414331e-8 k1=5.224851534e-01 lk1=-6.227372655e-9 k2=-7.144540537e-03 lk2=3.224478319e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.223655613e+00 ldsub=-4.419034005e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.205557218e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.404503811e-7 nfactor='7.798850790e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.101323326e-6 eta0=-7.462418332e-03 leta0=2.249307616e-7 etab=-1.632744345e+00 letab=7.978799692e-7 u0=1.148324636e-02 lu0=-2.564877967e-9 ua=-1.059609635e-10 lua=-5.351404061e-16 ub=4.864006036e-19 lub=3.665394455e-25 uc=-9.754060033e-11 luc=3.244585840e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.249860650e+04 lvsat=3.449316359e-2 a0=1.663177455e+00 la0=-4.477281531e-7 ags=-3.493192283e-01 lags=7.818591911e-07 pags=-1.776356839e-27 a1=0.0 a2=1.047418086e+00 la2=-4.690021102e-8 b0=-8.575503616e-17 lb0=8.480058261e-23 b1=-3.565229431e-20 lb1=3.525548427e-26 keta=1.023393023e-02 lketa=-2.366260124e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.536347840e+00 lpclm=-7.221227228e-7 pdiblc1=6.191336573e-02 lpdiblc1=-2.265833997e-8 pdiblc2=7.533057929e-04 lpdiblc2=-3.197073994e-10 pdiblcb=-1.477237207e-02 lpdiblcb=-1.011379443e-8 drout=1.036997061e+00 ldrout=-3.658528362e-8 pscbe1=8.230739141e+08 lpscbe1=-3.636238561e+1 pscbe2=3.809477986e-09 lpscbe2=5.307539814e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.632459620e+00 lbeta0=1.024241563e-6 agidl=2.197045537e-09 lagidl=-1.074069652e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.670956386e-01 lkt1=-1.183588529e-8 kt2=-6.206186670e-02 lkt2=1.335240081e-8 at=8.443425409e+04 lat=-2.242016604e-2 ute=-1.875821105e+00 lute=8.184494349e-7 ua1=-3.292299871e-09 lua1=2.830042980e-15 wua1=3.308722450e-30 pua1=3.308722450e-36 ub1=4.034982618e-18 lub1=-3.105147788e-24 wub1=6.162975822e-39 uc1=3.136276955e-10 luc1=-2.439630433e-16 puc1=2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.123 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.826083314e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.343176261e-8 k1=4.446623754e-01 lk1=3.181784882e-8 k2=1.132757422e-02 lk2=-5.805984424e-09 wk2=-2.081668171e-23 pk2=-9.540979118e-30 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.244403898e-01 ldsub=2.171402925e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-9.797583253e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.329269957e-7 nfactor='2.625212974e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.279129933e-7 eta0=4.169452362e-01 leta0=1.745059157e-8 etab=-1.210426333e-03 letab=2.719825911e-10 u0=4.591262030e-03 lu0=8.044064145e-10 ua=-1.330850367e-09 lua=6.367127645e-17 wua=-6.617444900e-30 ub=7.875179014e-19 lub=2.193322321e-25 uc=-6.000952568e-11 luc=1.409804193e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.833766079e+04 lvsat=-2.582274881e-3 a0=8.732071908e-01 la0=-6.153539006e-8 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=1.100021230e+00 la2=-7.261631000e-8 b0=1.715100723e-16 lb0=-4.096861098e-23 b1=7.130458861e-20 lb1=-1.703252708e-26 keta=-4.438001254e-02 lketa=3.036516966e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.930264200e-01 lpclm=2.699774716e-07 wpclm=-4.440892099e-22 ppclm=4.440892099e-28 pdiblc1=-3.561786926e-01 lpdiblc1=1.817343246e-07 wpdiblc1=-6.661338148e-22 ppdiblc1=-1.942890293e-28 pdiblc2=-8.000440691e-03 lpdiblc2=3.959736644e-09 ppdiblc2=-5.204170428e-30 pdiblcb=2.058549522e-01 lpdiblcb=-1.179718745e-7 drout=1.376341573e+00 ldrout=-2.024806355e-07 wdrout=-7.105427358e-21 pscbe1=6.996965507e+08 lpscbe1=2.395310605e+1 pscbe2=2.022856548e-08 lpscbe2=-2.719259489e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.553332902e+00 lbeta0=8.518424213e-8 agidl=0.0 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.663972928e-01 lkt1=1.344837144e-7 kt2=-1.748919269e-02 lkt2=-8.437842332e-9 at=1.056349506e+04 lat=1.369303193e-2 ute=4.030997005e-01 lute=-2.956465794e-07 pute=4.440892099e-28 ua1=4.600244176e-09 lua1=-1.028385029e-15 wua1=1.323488980e-29 ub1=-4.368480081e-18 lub1=1.003053022e-24 uc1=-2.690313562e-10 luc1=4.088148730e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.124 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.001582203e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.312662063e-8 k1=-7.003034297e-01 lk1=3.053158307e-7 k2=5.210617164e-01 lk2=-1.275661790e-07 pk2=1.110223025e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.906868453e+00 ldsub=-2.680784508e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.674043937e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.442801206e-8 nfactor='1.203208264e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.819105964e-06 wnfactor=5.684341886e-20 eta0=1.090917209e+00 leta0=-1.435410936e-7 etab=6.081955074e-02 letab=-1.454511803e-08 wetab=-8.500145032e-23 petab=1.669671346e-29 u0=1.672295362e-02 lu0=-2.093490755e-9 ua=7.735201398e-10 lua=-4.389997064e-16 ub=1.335696111e-18 lub=8.838890319e-26 uc=-1.074822148e-12 luc=2.030929986e-20 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.237216887e+05 lvsat=-1.103445762e-2 a0=-5.843766510e-01 la0=2.866376622e-7 ags=2.122259360e+00 lags=-1.472984366e-7 a1=0.0 a2=1.140496064e+00 la2=-8.228453375e-8 b0=0.0 b1=0.0 keta=-1.073852549e-01 lketa=1.808657922e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.739316293e-01 lpclm=-8.773797609e-9 pdiblc1=9.410904691e-01 lpdiblc1=-1.281443601e-7 pdiblc2=2.044747146e-02 lpdiblc2=-2.835616130e-9 pdiblcb=7.516267856e-02 lpdiblcb=-8.675341105e-8 drout=-6.083421165e-01 ldrout=2.716007575e-7 pscbe1=7.999088728e+08 lpscbe1=1.538866434e-2 pscbe2=1.279850067e-08 lpscbe2=-9.444399071e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025679629e+01 lbeta0=-3.217220576e-7 agidl=0.0 bgidl=1.818113540e+09 lbgidl=-1.381548261e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=4.646150296e-01 lkt1=-1.595681991e-7 kt2=4.349105275e-02 lkt2=-2.300419356e-8 at=1.364257274e+05 lat=-1.637167951e-2 ute=-2.646312955e+00 lute=4.327666216e-7 ua1=-7.134207826e-10 lua1=2.408901201e-16 ub1=4.952164236e-19 lub1=-1.587381621e-25 uc1=-2.797257078e-10 luc1=4.343604708e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.125 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.9e-07 wmax=8.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-6.678926379e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.963265331e-08 wvth0=-2.825746309e-07 pvth0=5.252214664e-14 k1=4.084085152e-01 lk1=1.299754278e-07 wk1=6.053131695e-07 pk1=-1.125095588e-13 k2=-3.370385465e-01 lk2=1.908693761e-08 wk2=3.965961450e-08 pk2=-7.371532548e-15 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.545913526e+00 ldsub=-4.138449893e-07 wdsub=-1.927334129e-06 pdsub=3.582335946e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.763281938e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.813951764e-08 wvoff=1.864483316e-07 pvoff=-3.465515139e-14 nfactor='-1.673535375e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.344769579e-06 wnfactor=1.598317132e-05 pnfactor=-2.970792053e-12 eta0=5.170531424e+00 leta0=-9.162691482e-07 weta0=-4.267190487e-06 peta0=7.931426957e-13 etab=4.499375087e-01 letab=-8.833471760e-08 wetab=-4.113870507e-07 petab=7.646451112e-14 u0=-3.699187191e-03 lu0=1.491622615e-09 wu0=7.596579014e-09 pu0=-1.411976141e-15 ua=-5.808584233e-09 lua=7.402223043e-16 wua=3.447316618e-15 pua=-6.407527398e-22 ub=5.914965134e-18 lub=-7.538617939e-25 wub=-3.510838116e-24 pub=6.525594806e-31 uc=-2.414450447e-10 luc=4.469996709e-17 wuc=2.081738630e-16 puc=-3.869327591e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.754167315e+05 lvsat=4.345557102e-02 wvsat=1.950249121e-01 pvsat=-3.624928042e-8 a0=-3.555136077e+00 la0=8.676682875e-07 wa0=4.040849822e-06 pa0=-7.510727564e-13 ags=1.250000055e+00 lags=-8.517666572e-15 a1=0.0 a2=2.507997991e+00 la2=-3.447456312e-07 wa2=-1.605527534e-06 pa2=2.984194027e-13 b0=0.0 b1=0.0 keta=-2.431940821e-01 lketa=4.515012654e-08 wketa=2.102704106e-07 pketa=-3.908296121e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.985881834e-01 lpclm=4.347037898e-09 wpclm=2.024469605e-08 ppclm=-3.762881655e-15 pdiblc1=3.539925496e+00 lpdiblc1=-6.240900108e-07 wpdiblc1=-2.906472543e-06 ppdiblc1=5.402260516e-13 pdiblc2=-4.333623387e-02 lpdiblc2=8.734402102e-09 wpdiblc2=4.067729445e-08 ppdiblc2=-7.560688720e-15 pdiblcb=-1.404858519e+01 lpdiblcb=2.529694214e-06 wpdiblcb=1.178113131e-05 ppdiblcb=-2.189758877e-12 drout=1.000000895e+00 ldrout=-1.395987859e-13 pscbe1=8.000000007e+08 lpscbe1=-1.075172424e-7 pscbe2=-3.264784285e-08 lpscbe2=7.407595996e-15 wpscbe2=3.449818553e-14 ppscbe2=-6.412177744e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.396250352e+00 lbeta0=-8.289871313e-09 wbeta0=-3.860875508e-08 pbeta0=7.176209307e-15 agidl=0.0 bgidl=1.000000270e+09 lbgidl=-4.199738693e-5 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.665503459e+00 lkt1=2.202933289e-07 wkt1=1.816984979e-06 pkt1=-3.377229981e-13 kt2=7.222637721e-01 lkt2=-1.514834916e-07 wkt2=-7.054793537e-07 pkt2=1.311274475e-13 at=-3.723674392e+05 lat=7.654958324e-02 wat=3.565018818e-01 pat=-6.626300477e-8 ute=-7.848584152e+00 lute=1.443279018e-06 wute=6.721547513e-06 pute=-1.249334036e-12 ua1=-6.341296857e-09 lua1=1.311193651e-15 wua1=6.106407618e-15 pua1=-1.134997984e-21 ub1=5.984608789e-18 lub1=-1.195031558e-24 wub1=-5.565425826e-24 pub1=1.034445698e-30 uc1=-1.544564348e-10 luc1=2.452491740e-17 wuc1=1.142158864e-16 puc1=-2.122930681e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.126 pmos lmin=2.0e-05 lmax=0.0001 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.127 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.110394410e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.886777775e-7 k1=4.210956021e-01 lk1=2.110826255e-7 k2=1.775005695e-02 lk2=2.994270855e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=5.082197684e-27 pcit=-2.710505431e-32 voff='-1.239825132e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.344269313e-6 nfactor='1.349753009e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.079466284e-5 eta0=0.08 etab=-0.07 u0=1.179712614e-02 lu0=-1.779861227e-8 ua=-8.962599665e-10 lua=1.912151425e-15 ub=1.670762721e-18 lub=-5.162101108e-24 uc=-1.282222813e-10 luc=4.509347416e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.679434284e+04 lvsat=1.066639228e+0 a0=1.542842824e+00 la0=-1.575978955e-6 ags=8.774092800e-02 lags=5.106970788e-7 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=-1.704051168e-07 lb0=1.361344325e-12 b1=-1.069304601e-10 lb1=8.542535445e-16 keta=4.015882949e-02 lketa=-3.357644528e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=1.914844237e-03 lpdiblc2=-1.274661131e-8 pdiblcb=-2.715221659e-01 lpdiblcb=9.299255256e-7 drout=0.56 pscbe1=8.000324548e+08 lpscbe1=-6.487344657e-1 pscbe2=1.314643402e-08 lpscbe2=-6.168183535e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.579227219e+01 lbeta0=-3.156696758e-4 agidl=-6.154969226e-08 lagidl=1.267496459e-12 wagidl=-5.293955920e-29 pagidl=-1.323488980e-33 bgidl=1000000000.0 cgidl=300.0 egidl=-4.229045954e-01 legidl=1.045227198e-05 pegidl=-7.105427358e-27 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.365713387e-01 lkt1=-3.355454267e-8 kt2=-6.266527973e-02 lkt2=8.233974711e-8 at=1.182508234e+05 lat=-9.446904559e-1 ute=-5.016829954e-02 lute=-6.558688149e-7 ua1=2.268269050e-09 lua1=-3.559399084e-15 ub1=-1.570431596e-18 lub1=6.826830664e-24 uc1=-4.378798232e-11 luc1=2.798238376e-16 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.128 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.067406195e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.525052071e-8 k1=4.556026508e-01 lk1=-6.458970099e-8 k2=1.888114602e-02 lk2=2.090658503e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.337794727e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.015363250e-7 nfactor='9.216209407e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-6.591748511e-6 eta0=0.08 etab=-0.07 u0=9.233736033e-03 lu0=2.679978022e-9 ua=-6.951832022e-10 lua=3.057752950e-16 ub=1.032606613e-18 lub=-6.395491904e-26 uc=-7.084610619e-11 luc=-7.436062681e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.668846287e+05 lvsat=-8.514108537e-1 a0=1.423035853e+00 la0=-6.188566371e-7 ags=1.271922909e-01 lags=1.955252693e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=-8.453595753e-04 lketa=-8.187316924e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.398542052e-01 lpclm=-7.900610979e-7 pdiblc1=0.39 pdiblc2=-1.382883923e-03 lpdiblc2=1.359851026e-8 pdiblcb=-2.485894473e-01 lpdiblcb=7.467190179e-7 drout=0.56 pscbe1=1.223533045e+09 lpscbe1=-3.383939895e+3 pscbe2=-1.692187543e-08 lpscbe2=1.785299800e-13 wpscbe2=-2.646977960e-29 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=3.454111638e+00 lbeta0=2.256438486e-5 agidl=1.929216340e-07 lagidl=-7.654418858e-13 bgidl=1000000000.0 cgidl=300.0 egidl=1.668713786e+00 legidl=-6.257395361e-06 pegidl=-1.421085472e-26 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.064088808e-01 lkt1=-2.745184978e-7 kt2=-4.842691408e-02 lkt2=-3.140870509e-8 at=-9.042369403e+04 lat=7.223831365e-1 ute=-1.644424595e-01 lute=2.570525935e-7 ua1=5.811130231e-10 lua1=9.919071081e-15 ub1=8.106627581e-19 lub1=-1.219542258e-23 pub1=-1.232595164e-44 uc1=-1.162365659e-11 luc1=2.286722078e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.129 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.059054255e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.193571586e-8 k1=4.427490850e-01 lk1=-1.331849770e-8 k2=2.173134058e-02 lk2=9.537529476e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.570387389e-01 ldsub=-1.184848914e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.130098824e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.186891293e-7 nfactor='8.071022804e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.023748026e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391144744e-01 letab=2.756886533e-7 u0=8.900325659e-03 lu0=4.009908663e-9 ua=-7.590571481e-10 lua=5.605601617e-16 ub=1.009458227e-18 lub=2.838098239e-26 uc=-7.555427377e-11 luc=1.134420574e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=53438.0 a0=1.240871201e+00 la0=1.077744766e-7 ags=7.206282245e-02 lags=4.154295521e-7 a1=0.0 a2=0.8 b0=0.0 b1=0.0 keta=6.416077653e-03 lketa=-3.715224604e-08 pketa=2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-5.457365877e-01 lpclm=2.343558448e-06 wpclm=-6.661338148e-22 ppclm=-2.220446049e-27 pdiblc1=0.39 pdiblc2=3.613575983e-03 lpdiblc2=-6.331718765e-9 pdiblcb=-9.757511029e-02 lpdiblcb=1.443424596e-7 drout=0.56 pscbe1=-3.954447050e+07 lpscbe1=1.654312115e+3 pscbe2=4.621586901e-08 lpscbe2=-7.331827470e-14 wpscbe2=1.058791184e-28 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.143313392e+01 lbeta0=-9.262897737e-6 agidl=1.380078841e-09 lagidl=-1.407522526e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.815048848e-01 lkt1=2.502969993e-08 wkt1=1.776356839e-21 kt2=-6.021807947e-02 lkt2=1.562472077e-08 wkt2=2.220446049e-22 at=1.020960915e+05 lat=-4.555326054e-2 ute=-1.321769333e-01 lute=1.283496039e-7 ua1=3.319292612e-09 lua1=-1.003171333e-15 ub1=-2.832123884e-18 lub1=2.335179770e-24 uc1=1.777277470e-11 luc1=-9.439132211e-17 wuc1=-2.584939414e-32 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.130 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.072527806e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.873285697e-8 k1=3.568093539e-01 lk1=1.576044552e-7 k2=5.659888429e-02 lk2=-5.980948219e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-2.484432034e-01 ldsub=1.013810956e-06 pdsub=1.776356839e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.430695179e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=7.958683643e-8 nfactor='8.417740844e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.713325134e-6 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=1.734723476e-22 peta0=-7.979727989e-29 etab=8.156999796e-01 letab=-1.623313170e-06 wetab=5.655198532e-22 petab=1.307981501e-27 u0=1.292093949e-02 lu0=-3.986569568e-9 ua=-3.091838044e-10 lua=-3.341794354e-16 ub=1.188535755e-18 lub=-3.277809421e-25 uc=-7.491430767e-11 luc=1.007139638e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.942857446e+04 lvsat=-1.191447383e-2 a0=1.378767846e+00 la0=-1.664840227e-7 ags=1.223252520e-01 lags=3.154641139e-7 a1=0.0 a2=6.022358887e-01 la2=3.933271080e-7 b0=0.0 b1=0.0 keta=-1.084892703e-02 lketa=-2.814396178e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=4.610337555e-01 lpclm=3.412231158e-7 pdiblc1=7.370933700e-01 lpdiblc1=-6.903235908e-7 pdiblc2=0.00043 pdiblcb=-0.025 drout=1.248972000e-01 ldrout=8.653629058e-7 pscbe1=7.981125877e+08 lpscbe1=-1.167887878e+1 pscbe2=9.524462383e-09 lpscbe2=-3.438368068e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=5.893237408e+00 lbeta0=1.755236233e-6 agidl=2.387521108e-10 lagidl=8.624279685e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.588881710e-01 lkt1=-1.995200383e-8 kt2=-5.612249362e-02 lkt2=7.479132955e-9 at=9.642825824e+04 lat=-3.428067692e-2 ute=9.019606480e-01 lute=-1.928415607e-06 wute=-8.881784197e-22 pute=4.440892099e-28 ua1=6.024083757e-09 lua1=-6.382649298e-15 ub1=-4.182471934e-18 lub1=5.020846495e-24 pub1=6.162975822e-45 uc1=-1.252175596e-10 luc1=1.899978642e-16 wuc1=2.067951531e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.131 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.056116434e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.250414331e-8 k1=5.224851534e-01 lk1=-6.227372655e-9 k2=-7.144540537e-03 lk2=3.224478319e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.223655613e+00 ldsub=-4.419034005e-07 wdsub=-3.552713679e-21 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.205557218e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.404503811e-7 nfactor='7.798850790e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.101323326e-06 wnfactor=2.842170943e-20 eta0=-7.462418332e-03 leta0=2.249307616e-7 etab=-1.632744345e+00 letab=7.978799692e-7 u0=1.148324636e-02 lu0=-2.564877967e-9 ua=-1.059609635e-10 lua=-5.351404061e-16 ub=4.864006036e-19 lub=3.665394455e-25 uc=-9.754060033e-11 luc=3.244585840e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.249860650e+04 lvsat=3.449316359e-2 a0=1.663177455e+00 la0=-4.477281531e-7 ags=-3.493192283e-01 lags=7.818591911e-07 pags=-8.881784197e-28 a1=0.0 a2=1.047418086e+00 la2=-4.690021102e-8 b0=-8.575503616e-17 lb0=8.480058261e-23 b1=-3.565229431e-20 lb1=3.525548427e-26 keta=1.023393023e-02 lketa=-2.366260124e-08 pketa=2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.536347840e+00 lpclm=-7.221227228e-7 pdiblc1=6.191336573e-02 lpdiblc1=-2.265833997e-8 pdiblc2=7.533057929e-04 lpdiblc2=-3.197073994e-10 pdiblcb=-1.477237207e-02 lpdiblcb=-1.011379443e-8 drout=1.036997061e+00 ldrout=-3.658528362e-8 pscbe1=8.230739141e+08 lpscbe1=-3.636238561e+1 pscbe2=3.809477986e-09 lpscbe2=5.307539814e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=6.632459620e+00 lbeta0=1.024241563e-6 agidl=2.197045537e-09 lagidl=-1.074069652e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.670956386e-01 lkt1=-1.183588529e-8 kt2=-6.206186670e-02 lkt2=1.335240081e-08 wkt2=-2.220446049e-22 at=8.443425409e+04 lat=-2.242016604e-2 ute=-1.875821105e+00 lute=8.184494349e-7 ua1=-3.292299871e-09 lua1=2.830042980e-15 wua1=-3.308722450e-30 pua1=-1.654361225e-36 ub1=4.034982618e-18 lub1=-3.105147788e-24 pub1=-3.081487911e-45 uc1=3.136276955e-10 luc1=-2.439630433e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.132 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.826083314e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.343176261e-8 k1=4.446623754e-01 lk1=3.181784882e-8 k2=1.132757422e-02 lk2=-5.805984424e-09 wk2=3.469446952e-24 pk2=-6.071532166e-30 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.244403898e-01 ldsub=2.171402925e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-9.797583253e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.329269957e-7 nfactor='2.625212974e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.279129933e-7 eta0=4.169452362e-01 leta0=1.745059157e-8 etab=-1.210426333e-03 letab=2.719825911e-10 u0=4.591262030e-03 lu0=8.044064145e-10 ua=-1.330850367e-09 lua=6.367127645e-17 ub=7.875179014e-19 lub=2.193322321e-25 uc=-6.000952568e-11 luc=1.409804193e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.833766079e+04 lvsat=-2.582274881e-3 a0=8.732071908e-01 la0=-6.153539006e-8 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=1.100021230e+00 la2=-7.261631000e-8 b0=1.715100723e-16 lb0=-4.096861098e-23 b1=7.130458861e-20 lb1=-1.703252708e-26 keta=-4.438001254e-02 lketa=3.036516966e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.930264200e-01 lpclm=2.699774716e-07 ppclm=-3.330669074e-28 pdiblc1=-3.561786926e-01 lpdiblc1=1.817343246e-07 wpdiblc1=-3.330669074e-22 ppdiblc1=1.387778781e-29 pdiblc2=-8.000440691e-03 lpdiblc2=3.959736644e-09 wpdiblc2=-4.336808690e-25 ppdiblc2=6.830473687e-30 pdiblcb=2.058549522e-01 lpdiblcb=-1.179718745e-07 ppdiblcb=5.551115123e-29 drout=1.376341573e+00 ldrout=-2.024806355e-7 pscbe1=6.996965507e+08 lpscbe1=2.395310605e+1 pscbe2=2.022856548e-08 lpscbe2=-2.719259489e-15 wpscbe2=-5.293955920e-29 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.553332902e+00 lbeta0=8.518424213e-8 agidl=0.0 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.663972928e-01 lkt1=1.344837144e-7 kt2=-1.748919269e-02 lkt2=-8.437842332e-9 at=1.056349506e+04 lat=1.369303193e-2 ute=4.030997005e-01 lute=-2.956465794e-7 ua1=4.600244176e-09 lua1=-1.028385029e-15 ub1=-4.368480081e-18 lub1=1.003053022e-24 uc1=-2.690313562e-10 luc1=4.088148730e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.133 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.001582203e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.312662063e-8 k1=-7.003034297e-01 lk1=3.053158307e-7 k2=5.210617164e-01 lk2=-1.275661790e-07 wk2=4.440892099e-22 pk2=-2.775557562e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.906868453e+00 ldsub=-2.680784508e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.674043937e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.442801206e-8 nfactor='1.203208264e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.819105964e-6 eta0=1.090917209e+00 leta0=-1.435410936e-07 weta0=3.552713679e-21 etab=6.081955074e-02 letab=-1.454511803e-08 wetab=-5.898059818e-23 petab=-1.138412281e-29 u0=1.672295362e-02 lu0=-2.093490755e-9 ua=7.735201398e-10 lua=-4.389997064e-16 ub=1.335696111e-18 lub=8.838890319e-26 uc=-1.074822148e-12 luc=2.030929986e-20 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.237216887e+05 lvsat=-1.103445762e-2 a0=-5.843766510e-01 la0=2.866376622e-7 ags=2.122259360e+00 lags=-1.472984366e-7 a1=0.0 a2=1.140496064e+00 la2=-8.228453375e-8 b0=0.0 b1=0.0 keta=-1.073852549e-01 lketa=1.808657922e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.739316293e-01 lpclm=-8.773797609e-9 pdiblc1=9.410904691e-01 lpdiblc1=-1.281443601e-7 pdiblc2=2.044747146e-02 lpdiblc2=-2.835616130e-9 pdiblcb=7.516267856e-02 lpdiblcb=-8.675341105e-8 drout=-6.083421165e-01 ldrout=2.716007575e-7 pscbe1=7.999088728e+08 lpscbe1=1.538866434e-2 pscbe2=1.279850067e-08 lpscbe2=-9.444399071e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025679629e+01 lbeta0=-3.217220576e-7 agidl=0.0 bgidl=1.818113540e+09 lbgidl=-1.381548261e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=4.646150296e-01 lkt1=-1.595681991e-07 pkt1=2.220446049e-28 kt2=4.349105275e-02 lkt2=-2.300419356e-8 at=1.364257274e+05 lat=-1.637167951e-2 ute=-2.646312955e+00 lute=4.327666216e-7 ua1=-7.134207826e-10 lua1=2.408901201e-16 pua1=4.135903063e-37 ub1=4.952164236e-19 lub1=-1.587381621e-25 pub1=-1.925929944e-46 uc1=-2.797257078e-10 luc1=4.343604708e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.134 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.5e-07 wmax=7.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-7.182488639e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.027294157e-08 wvth0=-2.404958605e-07 pvth0=4.470096560e-14 k1=4.032537413e-01 lk1=1.309335456e-07 wk1=6.096206119e-07 pk1=-1.133101831e-13 k2=-1.270326679e-01 lk2=-1.994685504e-08 wk2=-1.358259178e-07 pk2=2.524596334e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.562326471e+00 ldsub=-4.168956634e-07 wdsub=-1.941049147e-06 pdsub=3.607828049e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.087394108e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.345443390e-07 wvoff=5.299440526e-07 pvoff=-9.850070106e-14 nfactor='-1.687146450e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.370068486e-06 wnfactor=1.609690846e-05 pnfactor=-2.991932376e-12 eta0=5.170532605e+00 leta0=-9.162693676e-07 weta0=-4.267191473e-06 peta0=7.931428791e-13 etab=4.534408311e-01 letab=-8.898588015e-08 wetab=-4.143145040e-07 petab=7.700863687e-14 u0=-2.271727163e-03 lu0=1.226300619e-09 wu0=6.403762010e-09 pu0=-1.190267245e-15 ua=-5.808672994e-09 lua=7.402388024e-16 wua=3.447390789e-15 pua=-6.407665260e-22 ub=5.914943214e-18 lub=-7.538577197e-25 wub=-3.510819799e-24 pub=6.525560761e-31 uc=-2.432178282e-10 luc=4.502947436e-17 wuc=2.096552399e-16 puc=-3.896861943e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.916160934e+04 lvsat=2.184723147e-02 wvsat=9.787957447e-02 pvsat=-1.819287651e-8 a0=-3.555135937e+00 la0=8.676682617e-07 wa0=4.040849706e-06 pa0=-7.510727348e-13 ags=1.250000055e+00 lags=-8.517666572e-15 a1=0.0 a2=2.521670470e+00 la2=-3.472869348e-07 wa2=-1.616952558e-06 pa2=3.005429719e-13 b0=0.0 b1=0.0 keta=-2.431940735e-01 lketa=4.515012496e-08 wketa=2.102704034e-07 pketa=-3.908295989e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.984157820e-01 lpclm=4.379082144e-09 wpclm=2.038875844e-08 ppclm=-3.789658532e-15 pdiblc1=3.564676665e+00 lpdiblc1=-6.286905107e-07 wpdiblc1=-2.927155165e-06 ppdiblc1=5.440703305e-13 pdiblc2=-4.368263680e-02 lpdiblc2=8.798788014e-09 wpdiblc2=4.096675636e-08 ppdiblc2=-7.614491005e-15 pdiblcb=-1.414891189e+01 lpdiblcb=2.548341936e-06 wpdiblcb=1.186496650e-05 ppdiblcb=-2.205341324e-12 drout=1.000000895e+00 ldrout=-1.395988072e-13 wdrout=-8.526512829e-20 pdrout=1.421085472e-26 pscbe1=8.000000007e+08 lpscbe1=-1.075172424e-7 pscbe2=-3.294162523e-08 lpscbe2=7.462201327e-15 wpscbe2=3.474367655e-14 ppscbe2=-6.457807160e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.396579140e+00 lbeta0=-8.350983044e-09 wbeta0=-3.888349715e-08 pbeta0=7.227275615e-15 agidl=0.0 bgidl=1.000000270e+09 lbgidl=-4.199739456e-5 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-2.760146201e+00 lkt1=4.237545753e-07 wkt1=2.731692537e-06 pkt1=-5.077396918e-13 kt2=7.282715491e-01 lkt2=-1.526001571e-07 wkt2=-7.104995844e-07 pkt2=1.320605577e-13 at=-3.754033662e+05 lat=7.711387099e-02 wat=3.590387691e-01 pat=-6.673453602e-8 ute=-7.905824039e+00 lute=1.453918196e-06 wute=6.769378422e-06 pute=-1.258224367e-12 ua1=-6.393298287e-09 lua1=1.320859156e-15 wua1=6.149861156e-15 pua1=-1.143074693e-21 ub1=6.032003283e-18 lub1=-1.203840772e-24 wub1=-5.605029708e-24 pub1=1.041806872e-30 uc1=-1.554290835e-10 luc1=2.470570361e-17 wuc1=1.150286531e-16 puc1=-2.138037575e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.135 pmos lmin=2.0e-05 lmax=0.0001 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.136 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.136828158e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=9.170585294e-07 wvth0=2.103127143e-08 pvth0=-4.203913506e-13 k1=4.806021126e-01 lk1=-9.783852781e-07 wk1=-4.734468894e-08 pk1=9.463668324e-13 k2=-3.958080703e-02 lk2=1.175921896e-06 wk2=4.561369666e-08 pk2=-9.117662528e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=8.470329473e-28 pcit=-8.131516294e-32 voff='-1.894300151e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.742648538e-05 wvoff=5.207147233e-07 pvoff=-1.040849891e-11 nfactor='1.527600031e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.634427302e-05 wnfactor=-1.414990040e-06 pnfactor=2.828405196e-11 eta0=0.08 etab=-0.07 u0=1.629734614e-02 lu0=-1.077529249e-07 wu0=-3.580474042e-09 pu0=7.156963016e-14 ua=-7.744305291e-10 lua=-5.230813610e-16 wua=-9.693018063e-17 pua=1.937524780e-21 ub=1.229356260e-18 lub=3.661115263e-24 wub=3.511926915e-25 pub=-7.019945055e-30 uc=-4.796256430e-10 luc=7.475090855e-15 wuc=2.795842454e-16 puc=-5.588573135e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-9.584995976e+05 lvsat=2.076155172e+01 wvsat=7.839215355e-01 pvsat=-1.566970566e-5 a0=3.053401515e-01 la0=2.316030109e-05 wa0=9.845843511e-07 pa0=-1.968072860e-11 ags=-2.851467686e-01 lags=7.964300770e-06 wags=2.966776549e-07 pags=-5.930251076e-12 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=5.990387363e-07 lb0=-1.401896883e-11 wb0=-6.121864572e-13 pb0=1.223691551e-17 b1=1.703936494e-08 lb1=-3.418808162e-13 wb1=-1.364196984e-14 pb1=2.726875616e-19 keta=1.295143122e-01 lketa=-2.121879580e-06 wketa=-7.109318784e-08 pketa=1.421072490e-12 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 ppclm=1.332267630e-27 pdiblc1=0.39 pdiblc2=2.033233594e-03 lpdiblc2=-1.511308078e-08 wpdiblc2=-9.419317700e-11 ppdiblc2=1.882815170e-15 pdiblcb=-9.652811730e-01 lpdiblcb=1.479738413e-05 wpdiblcb=5.519699288e-07 ppdiblcb=-1.103325515e-11 drout=0.56 pscbe1=8.005164348e+08 lpscbe1=-1.032294826e+01 wpscbe1=-3.850651552e-01 ppscbe1=7.697017329e-6 pscbe2=7.697886426e-08 lpscbe2=-1.337619985e-12 wpscbe2=-5.078648581e-14 ppscbe2=1.015164463e-18 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=1.324310849e+01 lbeta0=3.349513260e-04 wbeta0=2.589683072e-05 pbeta0=-5.176483827e-10 agidl=-1.017691499e-06 lagidl=2.037969073e-11 wagidl=7.607274562e-13 pagidl=-1.520608223e-17 bgidl=1000000000.0 cgidl=300.0 egidl=-8.220688001e+00 legidl=1.663211508e-04 wegidl=6.204088029e-06 pegidl=-1.240127091e-10 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.203490209e-01 lkt1=-2.356707345e-06 wkt1=-9.246903295e-08 pkt1=1.848351479e-12 kt2=-2.494669610e-02 lkt2=-6.716121177e-07 wkt2=-3.000973495e-08 pkt2=5.998606906e-13 at=7.314087702e+05 lat=-1.320102494e+01 wat=-4.878419519e-01 pat=9.751409357e-6 ute=-9.142973343e+00 lute=1.810990291e-04 wute=7.234435734e-06 pute=-1.446081954e-10 ua1=-2.010032758e-08 lua1=4.435635709e-13 wua1=1.779694758e-14 pua1=-3.557408716e-19 ub1=1.442100735e-17 lub1=-3.128239635e-22 wub1=-1.272314063e-23 pub1=2.543212041e-28 uc1=7.075481051e-10 luc1=-1.473853554e-14 wuc1=-5.977795205e-16 puc1=1.194893712e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.137 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.046815447e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.979586828e-07 wvth0=-1.638245257e-08 pvth0=-1.214979733e-13 k1=3.847944230e-01 lk1=-2.129901005e-07 wk1=5.633658385e-08 pk1=1.180706227e-13 k2=7.103734872e-02 lk2=2.922078298e-07 wk2=-4.149662230e-08 pk2=-2.158532389e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='9.589002304e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-5.367361551e-06 wvoff=-1.346733211e-06 pvoff=4.510299866e-12 nfactor='9.080066650e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.684576446e-05 wnfactor=1.083181730e-07 pnfactor=1.611454067e-11 eta0=0.08 etab=-0.07 u0=1.548337290e-02 lu0=-1.012501985e-07 wu0=-4.972348583e-09 pu0=8.268913493e-14 ua=1.585742728e-09 lua=-1.937819869e-14 wua=-1.814754850e-15 pua=1.566100275e-20 ub=6.987221940e-19 lub=7.900281830e-24 wub=2.656457888e-25 pub=-6.336521971e-30 uc=4.684238456e-10 luc=-9.875326261e-17 wuc=-4.290550376e-16 puc=7.265397324e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.301030589e+06 lvsat=-1.326728120e+01 wvsat=-2.414033277e+00 pvsat=9.878339601e-6 a0=5.201663070e+00 la0=-1.595578619e-05 wa0=-3.006358944e-06 pa0=1.220239856e-11 ags=1.347436732e+00 lags=-5.078196578e-06 wags=-9.708533225e-07 pags=4.195889124e-12 a1=0.0 a2=0.8 b0=-8.636340129e-07 lb0=-2.333866379e-12 wb0=6.871262206e-13 pb0=1.856875437e-18 b1=1.949726913e-07 lb1=-1.763367029e-12 wb1=-1.551245626e-13 pb1=1.402973602e-18 keta=-1.258448413e-01 lketa=-8.184849989e-08 wketa=9.945233762e-08 pketa=5.860645772e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.873812691e+00 lpclm=-7.775450302e-05 wpclm=-7.664989318e-06 ppclm=6.123460321e-11 pdiblc1=0.39 pdiblc2=-2.547549491e-02 lpdiblc2=2.046505751e-07 wpdiblc2=1.916861134e-08 ppdiblc2=-1.520052259e-13 pdiblcb=-6.003656642e-01 lpdiblcb=1.188212157e-05 wpdiblcb=2.798808973e-07 ppdiblcb=-8.859571249e-12 drout=0.56 pscbe1=7.539444167e+09 lpscbe1=-5.384674054e+04 wpscbe1=-5.025077838e+03 ppscbe1=4.014931437e-2 pscbe2=-4.871533919e-07 lpscbe2=3.169159272e-12 wpscbe2=3.741265396e-13 ppscbe2=-2.379410459e-18 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-1.387094614e-09 lalpha0=1.188020555e-14 walpha0=1.183165191e-15 palpha0=-9.452152897e-21 alpha1=-1.387094614e-09 lalpha1=1.188020555e-14 walpha1=1.183165191e-15 palpha1=-9.452152897e-21 beta0=4.117415699e+02 lbeta0=-2.848601077e-03 wbeta0=-3.248424841e-04 pbeta0=2.284362407e-9 agidl=3.063395926e-06 lagidl=-1.222358617e-11 wagidl=-2.283812497e-12 pagidl=9.116351669e-18 bgidl=1000000000.0 cgidl=300.0 egidl=2.506206400e+01 legidl=-9.957042824e-05 wegidl=-1.861226409e-05 pegidl=7.424190184e-11 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-2.943739230e-01 lkt1=-2.564219025e-06 wkt1=-8.913747720e-08 pkt1=1.821736113e-12 kt2=-1.949679391e-01 lkt2=6.866654895e-07 wkt2=1.165912634e-07 pkt2=-5.713156268e-13 at=-1.776518596e+06 lat=6.834480753e+00 wat=1.341494198e+00 pat=-4.862919330e-6 ute=2.587998156e+01 lute=-9.869480461e-05 wute=-2.072151673e-05 pute=7.872827453e-11 ua1=5.314906596e-08 lua1=-1.416163116e-13 wua1=-4.182421985e-14 pua1=1.205648842e-19 ub1=-3.054091048e-17 lub1=4.637095299e-23 wub1=2.494400140e-23 pub1=-4.659669686e-29 uc1=-8.396166079e-09 luc1=5.798985360e-14 wuc1=6.670926411e-15 puc1=-4.611980963e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.138 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.929728280e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.681252418e-08 wvth0=-5.257583705e-08 pvth0=2.287273224e-14 k1=1.283183924e+00 lk1=-3.796549029e-06 wk1=-6.686684474e-07 pk1=3.010021442e-12 k2=-2.143982826e-01 lk2=1.430773456e-06 wk2=1.878699230e-07 pk2=-1.130766571e-12 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.377755770e-01 ldsub=-1.108010666e-06 wdsub=1.532619541e-08 pdsub=-6.113420107e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.807037659e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.750316414e-07 wvoff=-1.848278570e-07 pvoff=-1.243895421e-13 nfactor='3.988402289e-01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.782519177e-06 wnfactor=6.104157245e-06 pnfactor=-7.802081925e-12 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391329935e-01 letab=2.757625239e-07 wetab=1.473425771e-11 petab=-5.877303857e-17 u0=-2.685138258e-02 lu0=6.761763755e-08 wu0=2.844484561e-08 pu0=-5.060770848e-14 ua=-6.190868297e-09 lua=1.164169173e-14 wua=4.321668450e-15 pua=-8.816392061e-21 ub=2.570623141e-18 lub=4.335123017e-25 wub=-1.242097151e-24 pub=-3.223313906e-31 uc=7.864042300e-10 luc=-1.367135679e-15 wuc=-6.857931487e-16 puc=1.096748923e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.942369141e+05 lvsat=1.472660479e+00 wvsat=3.561800105e-01 pvsat=-1.171681076e-6 a0=-1.110743027e+00 la0=9.223581121e-06 wa0=1.870996016e-06 pa0=-7.252736314e-12 ags=1.749571257e+00 lags=-6.682258923e-06 wags=-1.334662616e-06 pags=5.647077100e-12 a1=0.0 a2=0.8 b0=-1.171699636e-06 lb0=-1.105032659e-12 wb0=9.322300075e-13 pb0=8.791882940e-19 b1=-4.081603290e-07 lb1=6.424521816e-13 wb1=3.247413373e-13 pb1=-5.111490896e-19 keta=-2.339630630e-01 lketa=3.494210314e-07 wketa=1.912509327e-07 pketa=-3.075662042e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-1.774215065e+01 lpclm=3.240198468e-05 wpclm=1.368184535e-05 ppclm=-2.391514520e-11 pdiblc1=0.39 pdiblc2=5.125638564e-02 lpdiblc2=-1.014229212e-07 wpdiblc2=-3.790566750e-08 ppdiblc2=7.565665270e-14 pdiblcb=4.768531366e+00 lpdiblcb=-9.533710729e-06 wpdiblcb=-3.871581367e-06 ppdiblcb=7.700072034e-12 drout=0.56 pscbe1=-1.255920101e+10 lpscbe1=2.632414227e+04 wpscbe1=9.960914179e+03 ppscbe1=-1.962785960e-2 pscbe2=6.053861159e-07 lpscbe2=-1.188838794e-12 wpscbe2=-4.448881502e-13 ppscbe2=8.875326668e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=3.074189227e-09 lalpha0=-5.915275728e-15 walpha0=-2.366330381e-15 palpha0=4.706323505e-21 alpha1=3.074189227e-09 lalpha1=-5.915275728e-15 walpha1=-2.366330381e-15 palpha1=4.706323505e-21 beta0=-6.277588731e+02 lbeta0=1.297831055e-03 wbeta0=5.085552230e-04 pbeta0=-1.039952705e-9 agidl=8.517741141e-09 lagidl=-3.807422157e-14 wagidl=-5.678881155e-15 pagidl=2.917283243e-20 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.164895998e+00 lkt1=9.081803661e-07 wkt1=5.437210046e-07 pkt1=-7.026540994e-13 kt2=-1.677425974e-02 lkt2=-2.412593213e-08 wkt2=-3.456485874e-08 pkt2=3.162649396e-14 at=-7.852348418e+05 lat=2.880378726e+00 wat=7.059800118e-01 pat=-2.327935859e-6 ute=-7.147168510e-01 lute=7.387990047e-06 wute=4.634815744e-07 pute=-5.775929648e-12 ua1=9.969868771e-09 lua1=3.061989271e-14 wua1=-5.291344705e-15 pua1=-2.516000546e-20 ub1=-1.685864092e-17 lub1=-8.205841577e-24 wub1=1.115980554e-23 pub1=8.386668487e-30 uc1=1.324591417e-08 luc1=-2.833759103e-14 wuc1=-1.052460031e-14 puc1=2.247091104e-20 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.139 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.458266875e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.105800686e-07 wvth0=-1.008061971e-07 pvth0=1.187966485e-13 k1=-1.875322662e+00 lk1=2.485309964e-06 wk1=1.775933339e-06 pk1=-1.851973712e-12 k2=9.789291513e-01 lk2=-9.425996770e-07 wk2=-7.338262517e-07 pk2=7.023673004e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-7.830572264e+00 ldsub=1.613220630e-05 wdsub=6.032508687e-06 pdsub=-1.202852794e-11 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.072526285e-02+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-5.596945040e-07 wvoff=-5.031070009e-07 pvoff=5.086262986e-13 nfactor='1.502724855e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.131148329e-05 wnfactor=-5.258669743e-06 pnfactor=1.479710379e-11 eta0=3.764988462e+00 leta0=-7.487078167e-06 weta0=-3.167805135e-06 peta0=6.300352600e-12 etab=1.297621799e+01 letab=-2.580896558e-05 wetab=-9.675175659e-06 petab=1.924263714e-11 u0=1.508548701e-02 lu0=-1.578934426e-08 wu0=-1.722161628e-09 pu0=9.390547209e-15 ua=-7.635836457e-10 lua=8.475281065e-16 wua=3.615305106e-16 pua=-9.401925179e-22 ub=6.477219506e-18 lub=-7.336200012e-24 wub=-4.207793143e-24 pub=5.576052397e-30 uc=5.727359548e-10 luc=-9.421772562e-16 wuc=-5.152847972e-16 puc=7.576299775e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.070857726e+05 lvsat=-7.177271727e-01 wvsat=-5.152903153e-01 pvsat=5.615601111e-7 a0=6.507966665e+00 la0=-5.929042025e-06 wa0=-4.080903423e-06 pa0=4.584817923e-12 ags=-1.826231482e+00 lags=4.295478703e-07 wags=1.550314605e-06 pags=-9.076754648e-14 a1=0.0 a2=-2.346909555e+00 la2=6.258794007e-06 wa2=2.346404996e-06 pa2=-4.666694505e-12 b0=-1.883178055e-06 lb0=3.100054259e-13 wb0=1.498297891e-12 pb0=-2.466471370e-19 b1=-1.477589475e-07 lb1=1.245476861e-13 wb1=1.175602694e-13 pb1=-9.909287907e-20 keta=8.430415854e-02 lketa=-2.835710976e-07 wketa=-7.570588825e-08 pketa=2.233762083e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.307511939e+00 lpclm=9.659974780e-06 wpclm=5.385203862e-06 ppclm=-7.414203836e-12 pdiblc1=5.829624753e+00 lpdiblc1=-1.081870648e-05 wpdiblc1=-4.051730004e-06 ppdiblc1=8.058364253e-12 pdiblc2=9.415235240e-05 lpdiblc2=3.321096633e-10 wpdiblc2=2.672077771e-10 ppdiblc2=-2.642337545e-16 pdiblcb=-2.974292909e+00 lpdiblcb=5.865760187e-06 wpdiblcb=2.346522322e-06 ppdiblcb=-4.666927852e-12 drout=-3.762780049e+00 ldrout=8.597447556e-06 wdrout=3.093121548e-06 pdrout=-6.151816653e-12 pscbe1=7.699666654e+08 lpscbe1=-1.858394578e+02 wpscbe1=2.239351502e+01 ppscbe1=1.385659882e-4 pscbe2=6.023023057e-09 lpscbe2=3.216480191e-15 wpscbe2=2.785822160e-15 ppscbe2=-2.832666530e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=2.406692809e+01 lbeta0=1.434273567e-06 wbeta0=-1.445938813e-05 pbeta0=2.553649582e-13 agidl=-1.138384321e-08 lagidl=1.507442503e-15 wagidl=9.247192538e-15 pagidl=-5.131877539e-22 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-9.349135889e-01 lkt1=4.507752512e-07 wkt1=3.787362950e-07 pkt1=-3.745209601e-13 kt2=-9.469036779e-03 lkt2=-3.865507092e-08 wkt2=-3.711851664e-08 pkt2=3.670538755e-14 at=1.110109726e+06 lat=-8.892152242e-01 wat=-8.065072765e-01 pat=6.802047344e-7 ute=7.003004925e+00 lute=-7.961555261e-06 wute=-4.854125050e-06 pute=4.800098638e-12 ua1=5.087427921e-08 lua1=-5.073366207e-14 wua1=-3.568380220e-14 pua1=3.528664149e-20 ub1=-4.321027080e-17 lub1=4.420412454e-23 wub1=3.105137539e-23 pub1=-3.117507805e-29 uc1=-2.059363702e-09 luc1=2.102616960e-15 wuc1=1.538849222e-15 puc1=-1.521721830e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.140 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.104160415e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.599140454e-08 wvth0=3.822484863e-08 pvth0=-1.868698175e-14 k1=7.633193985e-01 lk1=-1.239640101e-07 wk1=-1.916130238e-07 pk1=9.367385893e-14 k2=5.140453207e-02 lk2=-2.539840681e-08 wk2=-4.658293025e-08 pk2=2.277299711e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.646496638e+01 ldsub=-7.892922996e-06 wdsub=-1.212632216e-05 pdsub=5.928195113e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-4.485058758e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.267863893e-07 wvoff=2.223775740e-08 pvoff=-1.087137246e-14 nfactor='-1.632557774e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.692386050e-06 wnfactor=1.919392608e-05 pnfactor=-9.383334641e-12 eta0=-7.970553271e+00 leta0=4.117846987e-06 weta0=6.335610271e-06 peta0=-3.097289793e-12 etab=-2.595370628e+01 letab=1.268766863e-05 wetab=1.935029238e-05 petab=-9.459777436e-12 u0=-7.841390815e-03 lu0=6.882357411e-09 wu0=1.537510648e-08 pu0=-7.516428305e-15 ua=1.358769378e-09 lua=-1.251203128e-15 wua=-1.165371684e-15 pua=5.697152551e-22 ub=-3.070796135e-18 lub=2.105546215e-24 wub=2.830183984e-24 pub=-1.383592044e-30 uc=-7.211540753e-10 luc=3.373117779e-16 wuc=4.961606002e-16 puc=-2.425580326e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.182292441e+05 lvsat=9.840208790e-02 wvsat=1.040099539e-01 pvsat=-5.084734617e-8 a0=2.822831235e-01 la0=2.273496587e-07 wa0=1.098669910e-06 pa0=-5.371067587e-13 ags=-3.974890310e+00 lags=2.554292126e-06 wags=2.884584115e-06 pags=-1.410186636e-12 a1=0.0 a2=6.945708973e+00 la2=-2.930397677e-06 wa2=-4.692809993e-06 pa2=2.294174021e-12 b0=-3.104425716e-06 lb0=1.517660600e-12 wb0=2.469949397e-12 pb0=-1.207484162e-18 b1=-4.313340879e-08 lb1=2.108662955e-14 wb1=3.431788897e-14 pb1=-1.677698638e-20 keta=-3.630914091e-01 lketa=1.588449574e-07 wketa=2.970258531e-07 pketa=-1.452070288e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.787427606e+00 lpclm=-3.289218088e-06 wpclm=-4.177874586e-06 ppclm=2.042437549e-12 pdiblc1=-1.012314940e+01 lpdiblc1=4.956513295e-06 wpdiblc1=8.103460008e-06 ppdiblc1=-3.961538494e-12 pdiblc2=7.533057929e-04 lpdiblc2=-3.197073994e-10 pdiblcb=5.883813445e+00 lpdiblcb=-2.893755443e-06 wpdiblcb=-4.693044645e-06 ppdiblcb=2.294288736e-12 drout=8.812351559e+00 ldrout=-3.837722837e-06 wdrout=-6.186243096e-06 pdrout=3.024268662e-12 pscbe1=4.190874397e+08 lpscbe1=1.611344822e+02 wpscbe1=3.214205268e+02 ppscbe1=-1.571328529e-4 pscbe2=4.005175368e-09 lpscbe2=5.211869235e-15 wpscbe2=-1.557011422e-16 ppscbe2=7.611761738e-23 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.193336930e+01 lbeta0=-1.623331415e-05 wbeta0=-2.808618036e-05 pbeta0=1.373049099e-11 agidl=-1.949939707e-08 lagidl=9.532670247e-15 wagidl=1.726216706e-14 pagidl=-8.438955611e-21 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.670956386e-01 lkt1=-1.183588529e-8 kt2=-6.206186670e-02 lkt2=1.335240081e-8 at=3.793635449e+05 lat=-1.666022485e-01 wat=-2.346522322e-01 pat=1.147144368e-7 ute=-1.875821105e+00 lute=8.184494349e-7 ua1=-3.292299871e-09 lua1=2.830042980e-15 pua1=-2.481541838e-36 ub1=5.214699782e-18 lub1=-3.681876117e-24 wub1=-9.386089290e-25 pub1=4.588577471e-31 uc1=3.136276955e-10 luc1=-2.439630433e-16 puc1=2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.141 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.826083314e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.343176261e-8 k1=4.446623754e-01 lk1=3.181784882e-8 k2=1.132757422e-02 lk2=-5.805984424e-09 wk2=1.734723476e-24 pk2=4.336808690e-31 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.244403898e-01 ldsub=2.171402925e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-9.797583253e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.329269957e-7 nfactor='2.625212974e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.279129933e-7 eta0=4.169452362e-01 leta0=1.745059157e-8 etab=-1.210426333e-03 letab=2.719825911e-10 petab=-4.336808690e-31 u0=4.591262030e-03 lu0=8.044064145e-10 ua=-1.330850367e-09 lua=6.367127645e-17 ub=7.875179014e-19 lub=2.193322321e-25 uc=-6.000952568e-11 luc=1.409804193e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.833766079e+04 lvsat=-2.582274881e-3 a0=8.732071908e-01 la0=-6.153539006e-8 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=1.100021230e+00 la2=-7.261631000e-8 b0=1.715100723e-16 lb0=-4.096861098e-23 b1=7.130458861e-20 lb1=-1.703252708e-26 keta=-4.438001254e-02 lketa=3.036516966e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.930264200e-01 lpclm=2.699774716e-07 wpclm=-2.220446049e-22 ppclm=5.551115123e-29 pdiblc1=-3.561786926e-01 lpdiblc1=1.817343246e-07 wpdiblc1=-3.330669074e-22 ppdiblc1=2.081668171e-28 pdiblc2=-8.000440691e-03 lpdiblc2=3.959736644e-09 wpdiblc2=2.602085214e-24 ppdiblc2=1.951563910e-30 pdiblcb=2.058549522e-01 lpdiblcb=-1.179718745e-07 wpdiblcb=-2.220446049e-22 ppdiblcb=2.775557562e-29 drout=1.376341573e+00 ldrout=-2.024806355e-7 pscbe1=6.996965507e+08 lpscbe1=2.395310605e+1 pscbe2=2.022856548e-08 lpscbe2=-2.719259489e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.553332902e+00 lbeta0=8.518424213e-8 agidl=0.0 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.663972928e-01 lkt1=1.344837144e-7 kt2=-1.748919269e-02 lkt2=-8.437842332e-9 at=1.056349506e+04 lat=1.369303193e-2 ute=4.030997005e-01 lute=-2.956465794e-7 ua1=4.600244176e-09 lua1=-1.028385029e-15 ub1=-4.368480081e-18 lub1=1.003053022e-24 wub1=6.162975822e-39 uc1=-2.690313562e-10 luc1=4.088148730e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.142 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.209162380e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.068520287e-08 wvth0=2.458505071e-07 pvth0=-5.872631064e-14 k1=-1.995102558e+00 lk1=6.146044986e-07 wk1=1.030170672e-06 pk1=-2.460768685e-13 k2=1.394589345e+00 lk2=-3.362257236e-07 wk2=-6.949977990e-07 pk2=1.660141242e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=6.029553202e+00 ldsub=-1.252864157e-06 wdsub=-3.280098685e-06 pdsub=7.835171729e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='1.467241844e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.515879347e-07 wvoff=-1.618809309e-06 pvoff=3.866849796e-13 nfactor='3.392493300e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.048651128e-06 wnfactor=-1.741843339e-05 pnfactor=4.160741183e-12 eta0=1.005205903e+01 leta0=-2.284089039e-06 weta0=-7.129681574e-06 peta0=1.703067038e-12 etab=9.408004333e-01 letab=-2.247461515e-07 wetab=-7.001321498e-07 petab=1.672405666e-13 u0=3.110376392e-04 lu0=1.826823615e-09 wu0=1.305768141e-08 pu0=-3.119088359e-15 ua=-6.465954509e-09 lua=1.290293603e-15 wua=5.759885299e-15 pua=-1.375863801e-21 ub=8.708471314e-18 lub=-1.672745910e-24 wub=-5.865942153e-24 pub=1.401197602e-30 uc=-4.463702374e-10 luc=1.063880251e-16 wuc=3.542868288e-16 puc=-8.462849481e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.078596635e+04 lvsat=3.065018593e-02 wvsat=1.388421295e-01 pvsat=-3.316521947e-8 a0=-9.070193890e+00 la0=2.313644826e-06 wa0=6.751502883e-06 pa0=-1.612731494e-12 ags=2.122259350e+00 lags=-1.472984343e-07 wags=7.489404652e-15 pags=-1.788993842e-21 a1=0.0 a2=4.574808674e+00 la2=-9.026387868e-07 wa2=-2.732414667e-06 pa2=6.526918915e-13 b0=0.0 b1=0.0 keta=-5.489558726e-01 lketa=1.235645527e-07 wketa=3.513232980e-07 pketa=-8.392059619e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.306276543e-01 lpclm=1.570222884e-09 wpclm=3.445359515e-08 ppclm=-8.229930273e-15 pdiblc1=7.158198815e+00 lpdiblc1=-1.613225031e-06 wpdiblc1=-4.946468176e-06 ppdiblc1=1.181562853e-12 pdiblc2=-6.656347226e-02 lpdiblc2=1.794868799e-08 wpdiblc2=6.922782106e-08 ppdiblc2=-1.653644962e-14 pdiblcb=-2.512532612e+01 lpdiblcb=5.932887348e-06 wpdiblcb=2.005006330e-05 ppdiblcb=-4.789358620e-12 drout=-6.083463697e-01 ldrout=2.716017735e-07 wdrout=3.383973521e-12 pdrout=-8.083297542e-19 pscbe1=7.999088715e+08 lpscbe1=1.538896829e-02 wpscbe1=1.012386322e-06 ppscbe1=-2.418289185e-13 pscbe2=-6.099503773e-08 lpscbe2=1.668262261e-14 wpscbe2=5.871176260e-14 ppscbe2=-1.402447873e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.033939091e+01 lbeta0=-3.414514355e-07 wbeta0=-6.571410038e-08 pbeta0=1.569712716e-14 agidl=3.724644124e-08 lagidl=-8.897057420e-15 wagidl=-2.963408808e-14 pagidl=7.078694619e-21 bgidl=1.818113535e+09 lbgidl=-1.381548250e+02 wbgidl=3.757583618e-06 pbgidl=-8.975744247e-13 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-9.872052731e+00 lkt1=2.309551629e-06 wkt1=8.224080277e-06 pkt1=-1.964486056e-12 kt2=1.552549457e+00 lkt2=-3.834729746e-07 wkt2=-1.200640066e-06 pkt2=2.867968925e-13 at=-6.261514054e+05 lat=1.657851202e-01 wat=6.067231435e-01 pat=-1.449279573e-7 ute=-1.702407539e+01 lute=3.867182733e-06 wute=1.143926410e-05 pute=-2.732497016e-12 ua1=-1.377535434e-08 lua1=3.360994189e-15 wua1=1.039236170e-14 pua1=-2.482423440e-21 ub1=1.239997046e-17 lub1=-3.002426759e-24 wub1=-9.471684215e-24 pub1=2.262501209e-30 uc1=-5.240397428e-10 luc1=1.017953406e-16 wuc1=1.943816211e-16 puc1=-4.643193783e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.143 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-07 wmax=7.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='2.232296297e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.214577549e-07 wvth0=-9.895568626e-07 pvth0=1.649869292e-13 k1=3.720798198e+00 lk1=-3.859382602e-07 wk1=-2.029890744e-06 pk1=2.979243967e-13 k2=-2.409003659e+00 lk2=3.369005489e-07 wk2=1.679760406e-06 pk2=-2.586696819e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-8.000848692e+00 ldsub=1.228841869e-06 wdsub=6.463245402e-06 pdsub=-9.486021818e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.747618396e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.029847163e-06 wvoff=5.033343021e-06 pvoff=-8.108233243e-13 nfactor='-7.330312050e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.217224543e-05 wnfactor=6.099517547e-05 pnfactor=-9.995138001e-12 eta0=-1.784372389e+01 leta0=2.670962820e-06 weta0=1.404345731e-05 peta0=-2.060937969e-12 etab=-1.801253074e+00 letab=2.622943291e-07 wetab=1.379569570e-06 petab=-2.024776258e-13 u0=4.662702700e-02 lu0=-6.598024540e-09 wu0=-3.250116257e-08 pu0=5.034937987e-15 ua=1.278400471e-08 lua=-2.157803552e-15 wua=-1.134535263e-14 pua=1.664979728e-21 ub=-1.302000824e-17 lub=2.197532670e-24 wub=1.155424415e-23 pub=-1.695635049e-30 uc=8.977215665e-10 luc=-1.327283260e-16 wuc=-6.981012433e-16 puc=1.024593972e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.242060523e+05 lvsat=-5.455105230e-02 wvsat=-2.866983712e-01 pvsat=4.259127882e-8 a0=1.823837799e+01 la0=-2.529286762e-06 wa0=-1.329854943e-05 pa0=1.951619415e-12 ags=1.250000079e+00 lags=-1.228589142e-14 wags=-1.923450554e-14 pags=2.998081783e-21 a1=0.0 a2=-6.277752155e+00 la2=1.023658812e-06 wa2=5.384061670e-06 pa2=-7.902116248e-13 b0=0.0 b1=0.0 keta=8.908599478e-01 lketa=-1.316148749e-07 wketa=-6.920079252e-07 pketa=1.015551629e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=7.093695618e-01 lpclm=-1.290746246e-08 wpclm=-6.788850981e-08 ppclm=9.963896660e-15 pdiblc1=-1.236484697e+01 lpdiblc1=1.853121490e-06 wpdiblc1=9.746724286e-06 ppdiblc1=-1.430513897e-12 pdiblc2=1.792574833e-01 lpdiblc2=-2.593517378e-08 wpdiblc2=-1.364093079e-07 ppdiblc2=2.002061315e-14 pdiblcb=5.041997754e+01 lpdiblcb=-7.511459495e-06 wpdiblcb=-3.950746244e-05 ppdiblcb=5.798458010e-12 drout=1.000011818e+00 ldrout=-1.842213134e-12 wdrout=-8.690815633e-12 pdrout=1.354637433e-18 pscbe1=8.000000039e+08 lpscbe1=-6.168899536e-07 wpscbe1=-2.600036621e-06 ppscbe1=4.052677155e-13 pscbe2=1.561327559e-07 lpscbe2=-2.199549489e-14 wpscbe2=-1.156880607e-13 ppscbe2=1.697938402e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.184954496e+00 lbeta0=2.462003450e-08 wbeta0=1.294897247e-07 pbeta0=-1.900519131e-14 agidl=-9.565735425e-08 lagidl=1.491011181e-14 wagidl=7.610709551e-14 pagidl=-1.186281298e-20 bgidl=1.000000282e+09 lbgidl=-4.388798332e-05 wbgidl=-9.650329590e-06 pbgidl=1.504196167e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=2.282554161e+01 lkt1=-3.535449624e-06 wkt1=-1.762484357e-05 pkt1=2.642290272e-12 kt2=-3.138249688e+00 lkt2=4.498019627e-07 wkt2=2.365789776e-06 pkt2=-3.472238216e-13 at=1.578477725e+06 lat=-2.272998486e-01 wat=-1.195512013e+00 pat=1.754637164e-7 ute=2.893299129e+01 lute=-4.285551235e-06 wute=-2.254039350e-05 pute=3.308223781e-12 ua1=2.707408995e-08 lua1=-3.893343580e-15 wua1=-2.047752921e-14 pua1=3.005459716e-21 ub1=-2.447045059e-17 lub1=3.548426641e-24 wub1=1.866339365e-23 pub1=-2.739201632e-30 uc1=4.705542467e-10 luc1=-7.282219343e-17 wuc1=-3.830174561e-16 puc1=5.621496476e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.144 pmos lmin=2.0e-05 lmax=0.0001 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.145 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108621813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.532455644e-7 k1=4.171052081e-01 lk1=2.908460917e-7 k2=2.159455618e-02 lk2=-4.690448662e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=2.541098842e-27 pcit=2.710505431e-32 voff='-1.195937276e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.467000666e-6 nfactor='1.337826924e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.841077327e-5 eta0=0.08 etab=-0.07 u0=1.149534990e-02 lu0=-1.176644632e-8 ua=-9.044296180e-10 lua=2.075453526e-15 ub=1.700362603e-18 lub=-5.753769297e-24 uc=-1.046578370e-10 luc=-2.009187197e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.286628951e+04 lvsat=-2.540643246e-1 a0=1.625827411e+00 la0=-3.234747073e-6 ags=1.127460711e-01 lags=1.087252350e-8 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-06 wa2=1.776356839e-21 b0=-2.220025651e-07 lb0=2.392719013e-12 pb0=-1.694065895e-33 b1=-1.256728575e-09 lb1=2.383741859e-14 pb1=8.271806126e-37 keta=3.416681995e-02 lketa=-2.159909532e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 wpclm=-5.551115123e-23 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=1.906905271e-03 lpdiblc2=-1.258792035e-8 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=8.865952071e-09 lpscbe2=2.388016187e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.797495750e+01 lbeta0=-3.592990887e-4 agidl=2.567367474e-09 lagidl=-1.413111313e-14 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.443649873e-01 lkt1=1.222316870e-7 kt2=-6.519461656e-02 lkt2=1.328983321e-7 at=7.713361212e+04 lat=-1.228038641e-01 wat=-1.164153218e-16 ute=5.595779957e-01 lute=-1.284400824e-05 pute=3.552713679e-27 ua1=3.768264800e-09 lua1=-3.354261913e-14 wua1=-3.308722450e-30 pua1=2.646977960e-35 ub1=-2.642787222e-18 lub1=2.826200788e-23 uc1=-9.417115820e-11 luc1=1.286926591e-15 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.146 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.068786972e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.501020040e-8 k1=4.603509166e-01 lk1=-5.463825109e-8 k2=1.538364979e-02 lk2=2.713637080e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.472873697e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.816818865e-7 nfactor='9.225338883e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.233552538e-6 eta0=0.08 etab=-0.07 u0=8.814647214e-03 lu0=9.649338941e-9 ua=-8.481377777e-10 lua=1.625745332e-15 ub=1.054996270e-18 lub=-5.980215607e-25 uc=-1.070085284e-10 luc=-1.312504100e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.342054363e+04 lvsat=-1.882608877e-2 a0=1.169648264e+00 la0=4.096088288e-7 ags=4.536500838e-02 lags=5.491710742e-7 a1=0.0 a2=0.8 b0=5.791366221e-08 lb0=1.565046618e-13 b1=-1.307449963e-08 lb1=1.182480552e-13 wb1=3.308722450e-30 pb1=-6.617444900e-35 keta=7.536869066e-03 lketa=-3.247737421e-09 wketa=-1.387778781e-23 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.061808156e-01 lpclm=4.371028699e-06 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=2.327209668e-04 lpdiblc2=7.869204170e-10 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.461096001e-08 lpscbe2=-2.201595970e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.997217500e-10 lalpha0=-7.966640969e-16 alpha1=1.997217500e-10 lalpha1=-7.966640969e-16 beta0=-2.392487250e+01 lbeta0=2.150993062e-04 pbeta0=-2.842170943e-26 agidl=4.330612791e-10 lagidl=2.919581601e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.139217330e-01 lkt1=-1.209755144e-7 kt2=-3.860015032e-02 lkt2=-7.956140140e-8 at=2.264263863e+04 lat=3.125174394e-1 ute=-1.910932237e+00 lute=6.892576840e-6 ua1=-2.943994399e-09 lua1=2.008074701e-14 wua1=-1.654361225e-30 pua1=-6.617444900e-36 ub1=2.913039917e-18 lub1=-1.612277288e-23 uc1=5.506278879e-10 luc1=-3.864289165e-15 puc1=-2.481541838e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.147 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.063485550e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.386351842e-8 k1=3.863911154e-01 lk1=2.403777808e-7 k2=3.756574616e-02 lk2=-8.576786165e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.583304901e-01 ldsub=-1.190001542e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.285878909e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.082050964e-7 nfactor='8.585504846e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.681337744e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391132325e-01 letab=2.756836997e-7 u0=1.129776754e-02 lu0=-2.555052396e-10 ua=-3.948101738e-10 lua=-1.825195469e-16 ub=9.047694627e-19 lub=1.213642946e-27 uc=-1.333555795e-10 luc=1.037824576e-16 wuc=2.067951531e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.345823238e+04 lvsat=-9.875382428e-2 a0=1.398566000e+00 la0=-5.035142625e-7 ags=-4.042771799e-02 lags=8.913871067e-7 a1=0.0 a2=0.8 b0=7.857195977e-08 lb0=7.410139848e-14 b1=2.737045909e-08 lb1=-4.308162726e-14 keta=2.253544784e-02 lketa=-6.307511832e-08 pketa=2.775557562e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.074223900e-01 lpclm=3.278972801e-7 pdiblc1=0.39 pdiblc2=4.187393462e-04 lpdiblc2=4.491728403e-11 pdiblcb=-4.238870000e-01 lpdiblcb=7.933343877e-07 ppdiblcb=8.881784197e-28 drout=0.56 pscbe1=800000000.0 pscbe2=8.718970657e-09 lpscbe2=1.486419869e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-9.944350000e-11 lalpha0=3.966671938e-16 alpha1=-9.944350000e-11 lalpha1=3.966671938e-16 beta0=5.429614004e+01 lbeta0=-9.691414411e-5 agidl=9.014407177e-10 lagidl=1.051276909e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.356779703e-01 lkt1=-3.419271211e-8 kt2=-6.313133978e-02 lkt2=1.829032431e-8 at=1.615988244e+05 lat=-2.417607213e-1 ute=-9.311290905e-02 lute=-3.584681431e-7 ua1=2.873317563e-09 lua1=-3.123754152e-15 ub1=-1.891532201e-18 lub1=3.042040710e-24 wub1=-3.081487911e-39 uc1=-8.692813487e-10 luc1=1.799544192e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.148 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.081024143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.874549914e-8 k1=5.064919019e-01 lk1=1.512929702e-9 k2=-5.250837621e-03 lk2=-6.112426770e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.600000199e-01 ldsub=-1.966733887e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.854733267e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.224558331e-7 nfactor='7.974519768e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.466167851e-6 eta0=-4.835518650e-01 leta0=9.627162327e-07 weta0=4.180683577e-22 peta0=-7.372574773e-28 etab=2.386594872e-04 letab=-1.469097694e-9 u0=1.277578903e-02 lu0=-3.195097838e-9 ua=-2.787126111e-10 lua=-4.134225064e-16 ub=8.338866336e-19 lub=1.421903751e-25 uc=-1.183445084e-10 luc=7.392738859e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.599790864e+04 lvsat=3.541598979e-2 a0=1.034813481e+00 la0=2.199422095e-7 ags=2.529917783e-01 lags=3.078138731e-7 a1=0.0 a2=0.8 b0=1.262823559e-07 lb0=-2.078837708e-14 b1=9.908435342e-09 lb1=-8.351932082e-15 keta=-1.722971284e-02 lketa=1.601261680e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.149196182e-01 lpclm=-2.836747322e-7 pdiblc1=3.955978546e-01 lpdiblc1=-1.113340513e-8 pdiblc2=4.525213076e-04 lpdiblc2=-2.227064540e-11 pdiblcb=1.727740000e-01 lpdiblcb=-3.933467754e-7 drout=3.855974777e-01 ldrout=3.468639446e-7 pscbe1=800000000.0 pscbe2=9.759262277e-09 lpscbe2=-5.825849256e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.674544110e+00 lbeta0=1.776759381e-6 agidl=1.018141354e-09 lagidl=8.191745147e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.269668075e-01 lkt1=-5.151808255e-8 kt2=-5.925098613e-02 lkt2=1.057280534e-8 at=2.845269774e+04 lat=2.304961559e-2 ute=4.928361669e-01 lute=-1.523844682e-06 pute=8.881784197e-28 ua1=3.016514543e-09 lua1=-3.408554329e-15 ub1=-1.565341614e-18 lub1=2.393290035e-24 pub1=7.703719778e-46 uc1=4.482619664e-12 luc1=6.174124785e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.149 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.035203304e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.434645748e-09 wvth0=-1.319109069e-08 pvth0=1.304427385e-14 k1=-3.293797507e-01 lk1=8.280813307e-07 wk1=6.231275013e-07 pk1=-6.161920922e-13 k2=2.736935042e-01 lk2=-2.764509339e-07 wk2=-2.123264782e-07 pk2=2.099632845e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=7.802062121e+00 ldsub=-7.458118970e-06 wdsub=-5.667070156e-06 pdsub=5.603995665e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='1.635437654e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.172623408e-06 wvoff=-1.531596385e-06 pvoff=1.514549717e-12 nfactor='1.897092760e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.234018566e-05 wnfactor=-7.123924828e-06 pnfactor=7.044635545e-12 eta0=-4.439393457e+00 leta0=4.874529308e-06 weta0=3.702699827e-06 peta0=-3.661488778e-12 etab=-5.691544758e-03 letab=4.395103378e-09 wetab=2.881734220e-09 petab=-2.849660518e-15 u0=2.039780710e-01 lu0=-1.922692984e-07 wu0=-1.425621443e-07 pu0=1.409754276e-13 ua=2.666685468e-08 lua=-2.705908563e-14 wua=-2.003563686e-14 pua=1.981264022e-20 ub=7.139574768e-18 lub=-6.093315450e-24 wub=-4.782893190e-24 pub=4.729659589e-30 uc=-2.474564145e-10 luc=2.016022792e-16 wuc=1.429612030e-16 puc=-1.413700448e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.150047378e+05 lvsat=3.627345768e-01 wvsat=2.507300911e-01 pvsat=-2.479394652e-7 a0=5.855761333e+00 la0=-4.547348493e-06 wa0=-3.057038060e-06 pa0=3.023013226e-12 ags=-1.061952935e-01 lags=6.630031928e-07 wags=-4.920881480e-16 pags=4.866116399e-22 a1=0.0 a2=-4.480007950e+00 la2=5.221241461e-06 wa2=3.826455911e-06 pa2=-3.783867457e-12 b0=2.081769113e-07 lb0=-1.017714461e-13 wb0=7.306542202e-22 pb0=-7.225219627e-28 b1=2.892444750e-09 lb1=-1.414029464e-15 wb1=3.037671907e-25 pb1=-3.003856764e-31 keta=-2.464260546e-02 lketa=2.334300392e-08 wketa=4.467097925e-08 pketa=-4.417379126e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.354807759e+00 lpclm=-4.674146918e-06 wpclm=-3.109681710e-06 ppclm=3.075070953e-12 pdiblc1=1.351662203e+00 lpdiblc1=-9.565567569e-07 wpdiblc1=-4.524119689e-07 ppdiblc1=4.473766237e-13 pdiblc2=8.622179337e-03 lpdiblc2=-8.101000381e-09 wpdiblc2=-5.867205230e-09 ppdiblc2=5.801903235e-15 pdiblcb=-2.527982441e+00 lpdiblcb=2.277350246e-06 wpdiblcb=1.578975427e-06 ppdiblcb=-1.561401431e-12 drout=-4.514177379e+00 ldrout=5.192104307e-06 wdrout=3.750310063e-06 pdrout=-3.708569112e-12 pscbe1=-5.969729043e+09 lpscbe1=6.694381959e+03 wpscbe1=5.085062650e+03 ppscbe1=-5.028465903e-3 pscbe2=7.133571335e-07 lpscbe2=-6.963494119e-13 wpscbe2=-5.290641269e-13 ppscbe2=5.231756431e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.075903012e+00 lbeta0=5.335347604e-06 wbeta0=2.378045367e-06 pbeta0=-2.351577723e-12 agidl=2.425310328e-08 lagidl=-2.215718229e-14 wagidl=-1.536065976e-14 pagidl=1.518969562e-20 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.841236174e-01 lkt1=-9.388442793e-08 wkt1=-6.186576442e-08 pkt1=6.117719846e-14 kt2=-3.390872373e-01 lkt2=2.872944791e-07 wkt2=2.065562109e-07 pkt2=-2.042572403e-13 at=5.275063766e+05 lat=-4.704495958e-01 wat=-3.451107867e-01 pat=3.412697036e-7 ute=-2.288591904e+00 lute=1.226626094e-06 wute=3.077709884e-07 pute=-3.043454973e-13 ua1=-1.257732369e-08 lua1=1.201172448e-14 wua1=6.923118031e-15 pua1=-6.846063727e-21 ub1=2.015916203e-17 lub1=-1.908941988e-23 wub1=-1.208152876e-23 pub1=1.194706134e-29 uc1=1.632649380e-09 luc1=-1.548304017e-15 wuc1=-9.834915867e-16 puc1=9.725453254e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.150 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.017991114e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.979877251e-09 wvth0=2.638218138e-08 pvth0=-6.301911666e-15 k1=2.116092406e+00 lk1=-3.674366427e-07 wk1=-1.246255003e-06 pk1=2.976929325e-13 k2=-5.582008952e-01 lk2=1.302372811e-07 wk2=4.246529564e-07 pk2=-1.014368517e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.532536031e+01 ldsub=3.848184034e-06 wdsub=1.133414031e-05 pdsub=-2.707386096e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.087996508e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.114261850e-06 wvoff=3.063192770e-06 pvoff=-7.317048570e-13 nfactor='-1.648346362e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.992402570e-06 wnfactor=1.424784966e-05 pnfactor=-3.403383847e-12 eta0=1.034878691e+01 leta0=-2.354968430e-06 weta0=-7.405399655e-06 peta0=1.768927816e-12 etab=6.519319356e-03 letab=-1.574421762e-09 wetab=-5.763468440e-09 petab=1.376719706e-15 u0=-3.778066400e-01 lu0=9.214779328e-08 wu0=2.851242885e-07 pu0=-6.810763880e-14 ua=-5.507292573e-08 lua=1.290104082e-14 wua=4.007127372e-14 pua=-9.571825153e-21 ub=-1.204175267e-17 lub=3.283860093e-24 wub=9.565786380e-24 pub=-2.284979393e-30 uc=3.234587812e-10 luc=-7.750103253e-17 wuc=-2.859224059e-16 puc=6.829828510e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.608770739e+05 lvsat=-1.632317645e-01 wvsat=-5.014601823e-01 pvsat=1.197837937e-7 a0=-7.326760246e+00 la0=1.897190832e-06 wa0=6.114076120e-06 pa0=-1.460469363e-12 ags=1.005767372e+00 lags=1.193980046e-07 wags=9.841762960e-16 pags=-2.350910577e-22 a1=0.0 a2=1.136381686e+01 la2=-2.524329171e-06 wa2=-7.652911822e-06 pa2=1.828051047e-12 b0=2.131361386e-15 lb0=-5.091182942e-22 wb0=-1.461308256e-21 pb0=3.490627031e-28 b1=8.861044995e-19 lb1=-2.116637818e-25 wb1=-6.075327392e-25 pb1=1.451213454e-31 keta=7.544204007e-02 lketa=-2.558537674e-08 wketa=-8.934195851e-08 pketa=2.134111363e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-8.834201198e+00 lpclm=2.262433891e-06 wpclm=6.219363421e-06 ppclm=-1.485619340e-12 pdiblc1=-1.569694305e+00 lpdiblc1=4.716067989e-07 wpdiblc1=9.048239377e-07 ppdiblc1=-2.161352940e-13 pdiblc2=-2.373818778e-02 lpdiblc2=7.719012291e-09 wpdiblc2=1.173441046e-08 ppdiblc2=-2.802998626e-15 pdiblcb=4.441179090e+00 lpdiblcb=-1.129663751e-06 wpdiblcb=-3.157950854e-06 ppdiblcb=7.543397206e-13 drout=1.143588934e+01 ldrout=-2.605404811e-06 wdrout=-7.500620127e-06 pdrout=1.791673130e-12 pscbe1=1.433948360e+10 lpscbe1=-3.234182827e+03 wpscbe1=-1.017012530e+04 ppscbe1=2.429337831e-3 pscbe2=-1.398892992e-06 lpscbe2=3.362663069e-13 wpscbe2=1.058128254e-12 ppscbe2=-2.527550960e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.493202175e+01 lbeta0=-1.438493163e-06 wbeta0=-4.756090735e-06 pbeta0=1.136087394e-12 agidl=-4.120227075e-08 lagidl=9.841986413e-15 wagidl=3.072131952e-14 pagidl=-7.338401593e-21 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-9.323413352e-01 lkt1=1.741227678e-07 wkt1=1.237315288e-07 pkt1=-2.955575029e-14 kt2=5.365615486e-01 lkt2=-1.407839429e-07 wkt2=-4.131124218e-07 pkt2=9.868016420e-14 at=-9.151355499e+05 lat=2.348147628e-01 wat=6.902215733e-01 pat=-1.648732272e-7 ute=1.228641298e+00 lute=-4.928437007e-07 wute=-6.155419767e-07 pute=1.470345120e-13 ua1=2.317029182e-08 lua1=-5.464212308e-15 wua1=-1.384623606e-14 pua1=3.307450408e-21 ub1=-3.677505811e-17 lub1=8.744012315e-24 wub1=2.416305752e-23 pub1=-5.771829550e-30 uc1=-2.907074726e-09 luc1=6.710309070e-16 wuc1=1.966983173e-15 puc1=-4.698532706e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.151 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.794369863e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.807630180e-8 k1=-6.134766510e-01 lk1=2.845755181e-7 k2=4.624846070e-01 lk2=-1.135738648e-07 wk2=-1.110223025e-22 pk2=2.775557562e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.630409017e+00 ldsub=-2.020405853e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.038439192e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.701932152e-8 nfactor='1.056398954e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.468422564e-6 eta0=4.900000007e-01 leta0=-5.141975734e-17 etab=1.809698392e-03 letab=-4.494346021e-10 wetab=4.336808690e-25 petab=-1.626303259e-31 u0=1.782350564e-02 lu0=-2.356379616e-9 ua=1.258985607e-09 lua=-5.549628425e-16 ub=8.412917613e-19 lub=2.064872702e-25 uc=2.878584554e-11 luc=-7.112508390e-18 wuc=6.462348536e-33 puc=3.231174268e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.354238417e+05 lvsat=-1.382975091e-2 a0=-1.533380897e-02 la0=1.507103985e-7 ags=2.122259360e+00 lags=-1.472984367e-7 a1=0.0 a2=9.101975611e-01 la2=-2.727313031e-8 b0=0.0 b1=0.0 keta=-7.777436513e-02 lketa=1.101342597e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.768355118e-01 lpclm=-9.467448044e-9 pdiblc1=5.241829513e-01 lpdiblc1=-2.855766128e-8 pdiblc2=2.628226065e-02 lpdiblc2=-4.229372224e-09 wpdiblc2=2.775557562e-23 pdiblcb=1.765059758e+00 lpdiblcb=-4.904191263e-07 ppdiblcb=-4.440892099e-28 drout=-6.083418313e-01 ldrout=2.716006894e-7 pscbe1=7.999088729e+08 lpscbe1=1.538864396e-2 pscbe2=1.774695567e-08 lpscbe2=-2.126477355e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025125765e+01 lbeta0=-3.203990428e-7 agidl=-2.497675849e-09 lagidl=5.966198302e-16 bgidl=1.818113540e+09 lbgidl=-1.381548262e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.157772404e+00 lkt1=-3.251427011e-07 wkt1=8.881784197e-22 pkt1=1.110223025e-28 kt2=-5.770354749e-02 lkt2=1.168160598e-9 at=1.875627065e+05 lat=-2.858676971e-2 ute=-1.682167421e+00 lute=2.024611778e-7 ua1=1.624877580e-10 lua1=3.166184703e-17 ub1=-3.030938486e-19 lub1=3.195421259e-26 uc1=-2.633424711e-10 luc1=3.952258331e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.152 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=7.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.092643848e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.280651478e-09 wvth0=-8.412648320e-09 pvth0=1.563658943e-15 k1=1.606404155e-01 lk1=1.693383555e-07 wk1=6.246412223e-07 pk1=-1.161020640e-13 k2=4.596853226e-01 lk2=-1.244869467e-07 wk2=-4.591972097e-07 pk2=8.535098538e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.334815479e+00 ldsub=-5.391778692e-07 wdsub=-1.988875188e-06 pdsub=3.696722312e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='3.543980787e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.157770783e-07 wvoff=-2.640299745e-06 pvoff=4.907525136e-13 nfactor='8.429555484e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.532073346e-05 wnfactor=-5.651386404e-05 pnfactor=1.050423191e-11 eta0=6.713823862e+00 leta0=-1.156822141e-06 weta0=-4.267190562e-06 peta0=7.931427097e-13 etab=6.183274690e-01 letab=-1.150868368e-07 wetab=-4.245229134e-07 petab=7.890607392e-14 u0=-6.469423048e-03 lu0=1.921732297e-09 wu0=7.088718704e-09 pu0=-1.317580145e-15 ua=-7.055403364e-09 lua=9.345649958e-16 wua=3.447346496e-15 pua=-6.407582933e-22 ub=7.184684656e-18 lub=-9.517722683e-25 wub=-3.510819380e-24 pub=6.525559982e-31 uc=-3.266551770e-10 luc=5.823730427e-17 wuc=2.148209930e-16 puc=-3.992877797e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.183496227e+05 lvsat=3.194689359e-02 wvsat=1.178430763e-01 pvsat=-2.190349258e-8 a0=-5.016567780e+00 la0=1.095461645e-06 wa0=4.040849743e-06 pa0=-7.510727417e-13 ags=1.250000052e+00 lags=-8.145683239e-15 wags=4.785505325e-16 pags=-8.894573966e-23 a1=0.0 a2=3.165175715e+00 la2=-4.491514827e-07 wa2=-1.656793094e-06 pa2=3.079481325e-13 b0=0.0 b1=0.0 keta=-3.192415940e-01 lketa=5.700365207e-08 wketa=2.102704067e-07 pketa=-3.908296049e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.903016768e-01 lpclm=5.663515886e-09 wpclm=2.089112475e-08 ppclm=-3.883033357e-15 pdiblc1=4.729608978e+00 lpdiblc1=-8.130950725e-07 wpdiblc1=-2.999278144e-06 ppdiblc1=5.574758287e-13 pdiblc2=-5.998633668e-02 lpdiblc2=1.137960464e-08 wpdiblc2=4.197614767e-08 ppdiblc2=-7.802106568e-15 pdiblcb=-1.887086035e+01 lpdiblcb=3.295809265e-06 wpdiblcb=1.215731069e-05 ppdiblcb=-2.259679337e-12 drout=1.000000188e+00 ldrout=-3.018088357e-14 wdrout=-1.907957881e-14 pdrout=3.546320571e-21 pscbe1=8.000000016e+08 lpscbe1=-2.826652527e-07 wpscbe1=-8.396453857e-07 ppscbe1=1.560640335e-13 pscbe2=-4.676870923e-08 lpscbe2=9.650978605e-15 wpscbe2=3.559973552e-14 ppscbe2=-6.616922840e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=8.412055214e+00 lbeta0=-1.080078633e-08 wbeta0=-3.984156649e-08 pbeta0=7.405351963e-15 agidl=6.788365232e-08 lagidl=-1.242509642e-14 wagidl=-4.583267689e-14 pagidl=8.518919654e-21 bgidl=1.000000253e+09 lbgidl=-3.883447075e-05 wbgidl=1.217955780e-05 pbgidl=-2.263813972e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.321894018e+00 lkt1=1.030210562e-07 wkt1=3.800156765e-07 pkt1=-7.063351378e-14 kt2=1.011031791e+00 lkt2=-1.973600790e-07 wkt2=-7.280057794e-07 pkt2=1.353144342e-13 at=-5.182914647e+05 lat=9.973253917e-02 wat=3.678852243e-01 pat=-6.837882665e-8 ute=-1.059986113e+01 lute=1.880374504e-06 wute=6.936170982e-06 pute=-1.289226100e-12 ua1=-8.840781778e-09 lua1=1.708286927e-15 wua1=6.301389280e-15 pua1=-1.171239225e-21 ub1=8.262659774e-18 lub1=-1.556945610e-24 wub1=-5.743133568e-24 pub1=1.067476236e-30 uc1=-2.012074926e-10 luc1=3.195225987e-17 wuc1=1.178628755e-16 puc1=-2.190717267e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.153 pmos lmin=2.0e-05 lmax=0.0001 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.154 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108621813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.532455644e-7 k1=4.171052081e-01 lk1=2.908460917e-7 k2=2.159455618e-02 lk2=-4.690448662e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=-2.032879073e-26 pcit=-1.084202172e-31 voff='-1.195937276e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.467000666e-6 nfactor='1.337826924e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.841077327e-5 eta0=0.08 etab=-0.07 u0=1.149534990e-02 lu0=-1.176644632e-8 ua=-9.044296180e-10 lua=2.075453526e-15 ub=1.700362603e-18 lub=-5.753769297e-24 uc=-1.046578370e-10 luc=-2.009187197e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.286628951e+04 lvsat=-2.540643246e-1 a0=1.625827411e+00 la0=-3.234747073e-6 ags=1.127460711e-01 lags=1.087252350e-8 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=-2.220025651e-07 lb0=2.392719013e-12 b1=-1.256728575e-09 lb1=2.383741859e-14 wb1=2.481541838e-30 pb1=-1.985233470e-35 keta=3.416681995e-02 lketa=-2.159909532e-07 pketa=-1.776356839e-27 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=1.906905271e-03 lpdiblc2=-1.258792035e-08 wpdiblc2=-1.387778781e-23 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=8.865952071e-09 lpscbe2=2.388016187e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.797495750e+01 lbeta0=-3.592990887e-4 agidl=2.567367474e-09 lagidl=-1.413111313e-14 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.443649873e-01 lkt1=1.222316870e-7 kt2=-6.519461656e-02 lkt2=1.328983321e-7 at=7.713361212e+04 lat=-1.228038641e-1 ute=5.595779957e-01 lute=-1.284400824e-05 wute=8.881784197e-22 pute=-5.684341886e-26 ua1=3.768264800e-09 lua1=-3.354261913e-14 pua1=-2.117582368e-34 ub1=-2.642787222e-18 lub1=2.826200788e-23 pub1=9.860761315e-44 uc1=-9.417115820e-11 luc1=1.286926591e-15 puc1=-6.617444900e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.155 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.068786972e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.501020040e-8 k1=4.603509166e-01 lk1=-5.463825109e-8 k2=1.538364979e-02 lk2=2.713637080e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.472873697e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.816818865e-7 nfactor='9.225338883e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.233552538e-6 eta0=0.08 etab=-0.07 u0=8.814647214e-03 lu0=9.649338941e-9 ua=-8.481377777e-10 lua=1.625745332e-15 ub=1.054996270e-18 lub=-5.980215607e-25 uc=-1.070085284e-10 luc=-1.312504100e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.342054363e+04 lvsat=-1.882608877e-2 a0=1.169648264e+00 la0=4.096088288e-7 ags=4.536500838e-02 lags=5.491710742e-7 a1=0.0 a2=0.8 b0=5.791366221e-08 lb0=1.565046618e-13 b1=-1.307449963e-08 lb1=1.182480552e-13 pb1=2.117582368e-34 keta=7.536869066e-03 lketa=-3.247737421e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.061808156e-01 lpclm=4.371028699e-06 ppclm=-7.105427358e-27 pdiblc1=0.39 pdiblc2=2.327209668e-04 lpdiblc2=7.869204170e-10 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.461096001e-08 lpscbe2=-2.201595970e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.997217500e-10 lalpha0=-7.966640969e-16 alpha1=1.997217500e-10 lalpha1=-7.966640969e-16 beta0=-2.392487250e+01 lbeta0=2.150993062e-04 wbeta0=-5.684341886e-20 pbeta0=-6.821210263e-25 agidl=4.330612791e-10 lagidl=2.919581601e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.139217330e-01 lkt1=-1.209755144e-7 kt2=-3.860015032e-02 lkt2=-7.956140140e-8 at=2.264263863e+04 lat=3.125174394e-1 ute=-1.910932237e+00 lute=6.892576840e-6 ua1=-2.943994399e-09 lua1=2.008074701e-14 wua1=-1.323488980e-29 pua1=5.293955920e-35 ub1=2.913039917e-18 lub1=-1.612277288e-23 wub1=1.232595164e-38 pub1=-4.930380658e-44 uc1=5.506278879e-10 luc1=-3.864289165e-15 wuc1=-8.271806126e-31 puc1=-6.617444900e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.156 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.063485550e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.386351842e-8 k1=3.863911154e-01 lk1=2.403777808e-7 k2=3.756574616e-02 lk2=-8.576786165e-08 pk2=-4.440892099e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.583304901e-01 ldsub=-1.190001542e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.285878909e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.082050964e-07 wvoff=7.105427358e-21 nfactor='8.585504846e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.681337744e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391132325e-01 letab=2.756836997e-7 u0=1.129776754e-02 lu0=-2.555052396e-10 ua=-3.948101738e-10 lua=-1.825195469e-16 ub=9.047694627e-19 lub=1.213642946e-27 uc=-1.333555795e-10 luc=1.037824576e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.345823238e+04 lvsat=-9.875382428e-2 a0=1.398566000e+00 la0=-5.035142625e-7 ags=-4.042771799e-02 lags=8.913871067e-7 a1=0.0 a2=0.8 b0=7.857195977e-08 lb0=7.410139848e-14 b1=2.737045909e-08 lb1=-4.308162726e-14 keta=2.253544784e-02 lketa=-6.307511832e-08 wketa=1.110223025e-22 pketa=2.220446049e-28 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.074223900e-01 lpclm=3.278972801e-7 pdiblc1=0.39 pdiblc2=4.187393462e-04 lpdiblc2=4.491728403e-11 pdiblcb=-4.238870000e-01 lpdiblcb=7.933343877e-7 drout=0.56 pscbe1=800000000.0 pscbe2=8.718970657e-09 lpscbe2=1.486419869e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-9.944350000e-11 lalpha0=3.966671938e-16 alpha1=-9.944350000e-11 lalpha1=3.966671938e-16 beta0=5.429614004e+01 lbeta0=-9.691414411e-5 agidl=9.014407177e-10 lagidl=1.051276909e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.356779703e-01 lkt1=-3.419271211e-8 kt2=-6.313133979e-02 lkt2=1.829032431e-8 at=1.615988244e+05 lat=-2.417607213e-1 ute=-9.311290905e-02 lute=-3.584681431e-7 ua1=2.873317563e-09 lua1=-3.123754152e-15 ub1=-1.891532202e-18 lub1=3.042040710e-24 uc1=-8.692813487e-10 luc1=1.799544192e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.157 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.081024143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.874549914e-8 k1=5.064919019e-01 lk1=1.512929702e-9 k2=-5.250837621e-03 lk2=-6.112426770e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.600000199e-01 ldsub=-1.966733976e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.854733267e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.224558331e-7 nfactor='7.974519768e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.466167851e-6 eta0=-4.835518650e-01 leta0=9.627162327e-07 weta0=6.383782392e-22 peta0=-1.991462550e-27 etab=2.386594872e-04 letab=-1.469097694e-09 petab=6.938893904e-30 u0=1.277578903e-02 lu0=-3.195097838e-9 ua=-2.787126111e-10 lua=-4.134225064e-16 ub=8.338866336e-19 lub=1.421903751e-25 uc=-1.183445084e-10 luc=7.392738859e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.599790864e+04 lvsat=3.541598979e-2 a0=1.034813481e+00 la0=2.199422095e-7 ags=2.529917783e-01 lags=3.078138731e-7 a1=0.0 a2=0.8 b0=1.262823559e-07 lb0=-2.078837708e-14 b1=9.908435342e-09 lb1=-8.351932082e-15 keta=-1.722971284e-02 lketa=1.601261680e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.149196182e-01 lpclm=-2.836747322e-7 pdiblc1=3.955978546e-01 lpdiblc1=-1.113340513e-8 pdiblc2=4.525213076e-04 lpdiblc2=-2.227064540e-11 pdiblcb=1.727740000e-01 lpdiblcb=-3.933467754e-7 drout=3.855974777e-01 ldrout=3.468639446e-7 pscbe1=800000000.0 pscbe2=9.759262277e-09 lpscbe2=-5.825849256e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.674544110e+00 lbeta0=1.776759381e-6 agidl=1.018141354e-09 lagidl=8.191745147e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.269668075e-01 lkt1=-5.151808255e-8 kt2=-5.925098613e-02 lkt2=1.057280534e-8 at=2.845269774e+04 lat=2.304961559e-2 ute=4.928361669e-01 lute=-1.523844682e-06 pute=-3.552713679e-27 ua1=3.016514543e-09 lua1=-3.408554329e-15 ub1=-1.565341614e-18 lub1=2.393290035e-24 uc1=4.482619664e-12 luc1=6.174124785e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.158 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.054442900e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.246010562e-8 k1=5.794701714e-01 lk1=-7.065309168e-8 k2=-3.599095491e-02 lk2=2.978673710e-08 wk2=-1.110223025e-22 pk2=-5.551115123e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.635276000e-01 ldsub=7.154747378e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.984410505e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.639222613e-8 nfactor='8.580472176e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.065376009e-6 eta0=9.611039418e-01 leta0=-4.658605549e-7 etab=-1.488450021e-03 letab=2.387890846e-10 u0=-3.953040131e-03 lu0=1.334753945e-8 ua=-2.555715282e-09 lua=1.838237125e-15 ub=1.635833473e-19 lub=8.050331859e-25 uc=-3.894326448e-11 luc=-4.590119479e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.069252850e+04 lvsat=1.107521054e-3 a0=1.396980751e+00 la0=-1.381941390e-7 ags=-1.061952942e-01 lags=6.630031935e-7 a1=0.0 a2=1.100991363e+00 la2=-2.976413294e-7 b0=2.081769124e-07 lb0=-1.017714472e-13 b1=2.892444750e-09 lb1=-1.414029465e-15 keta=4.051134126e-02 lketa=-4.108577937e-08 wketa=8.326672685e-23 pketa=1.387778781e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=8.192448538e-01 lpclm=-1.890648279e-7 pdiblc1=6.918059423e-01 lpdiblc1=-3.040446968e-07 wpdiblc1=7.105427358e-21 pdiblc2=6.468668115e-05 lpdiblc2=3.612473816e-10 pdiblcb=-0.225 drout=9.557609593e-01 ldrout=-2.169536175e-7 pscbe1=1.446985488e+09 lpscbe1=-6.397845396e+2 pscbe2=-5.829857018e-08 lpscbe2=6.671776386e-14 ppscbe2=-1.588186776e-34 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.544352635e+00 lbeta0=1.905501825e-6 agidl=1.849125933e-09 lagidl=-2.561206190e-18 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.743566677e-01 lkt1=-4.655671468e-9 kt2=-3.781888407e-02 lkt2=-1.062075742e-8 at=2.415206960e+04 lat=2.730237773e-2 ute=-1.839698799e+00 lute=7.827291698e-7 ua1=-2.479750931e-09 lua1=2.026537710e-15 pua1=6.617444900e-36 ub1=2.537894393e-18 lub1=-1.664276955e-24 pub1=-6.162975822e-45 uc1=1.981977632e-10 luc1=-1.298178461e-16 wuc1=-8.271806126e-31 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.159 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.795119211e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.417140212e-8 k1=2.983925622e-01 lk1=6.675731910e-8 k2=6.116802299e-02 lk2=-1.771137242e-08 pk2=-1.110223025e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.205819134e+00 ldsub=-1.006188000e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.202390991e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.704863814e-8 nfactor='4.297447230e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.846639641e-8 eta0=-4.522078841e-01 leta0=2.250651974e-07 weta0=3.330669074e-22 peta0=-8.326672685e-29 etab=-1.886870119e-03 letab=4.335647182e-10 u0=3.805558220e-02 lu0=-7.189215745e-9 ua=3.372214182e-09 lua=-1.059749752e-15 wua=-1.323488980e-29 pua=-3.308722450e-36 ub=1.910230175e-18 lub=-4.885004854e-26 uc=-9.356751888e-11 luc=2.211403977e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.948254123e+04 lvsat=1.147644753e-2 a0=1.590800918e+00 la0=-2.329470036e-7 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=2.018182291e-01 la2=1.419374407e-7 b0=0.0 b1=0.0 keta=-5.486585336e-02 lketa=5.541269763e-09 wketa=4.440892099e-22 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.369246124e-01 lpclm=9.561406851e-8 pdiblc1=-2.499817842e-01 lpdiblc1=1.563670691e-07 ppdiblc1=-4.440892099e-28 pdiblc2=-6.623202468e-03 lpdiblc2=3.630755750e-09 wpdiblc2=-1.387778781e-23 pdiblcb=-1.647857919e-01 lpdiblcb=-2.943691991e-8 drout=4.960126660e-01 ldrout=7.803530650e-9 pscbe1=-4.939454606e+08 lpscbe1=3.090783733e+02 ppscbe1=-4.768371582e-19 pscbe2=1.444184156e-07 lpscbe2=-3.238448899e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=7.995122502e+00 lbeta0=2.185239603e-7 agidl=3.605683955e-09 lagidl=-8.612897264e-16 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.518752346e-01 lkt1=1.310148304e-7 kt2=-6.597515796e-02 lkt2=3.144000191e-9 at=9.157306403e+04 lat=-5.657723812e-3 ute=3.308550878e-01 lute=-2.783895088e-7 ua1=2.975146297e-09 lua1=-6.401978981e-16 ub1=-1.532522831e-18 lub1=3.256279136e-25 pub1=3.081487911e-45 uc1=-3.817149149e-11 luc1=-1.426400859e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.160 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.794369863e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.807630180e-8 k1=-6.134766510e-01 lk1=2.845755181e-7 k2=4.624846070e-01 lk2=-1.135738648e-07 wk2=-4.440892099e-22 pk2=1.110223025e-28 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.630409017e+00 ldsub=-2.020405853e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.038439192e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.701932152e-8 nfactor='1.056398954e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.468422564e-6 eta0=4.900000007e-01 leta0=-5.142197779e-17 etab=1.809698392e-03 letab=-4.494346021e-10 wetab=-3.469446952e-24 petab=-4.336808690e-31 u0=1.782350564e-02 lu0=-2.356379616e-9 ua=1.258985607e-09 lua=-5.549628425e-16 ub=8.412917613e-19 lub=2.064872702e-25 uc=2.878584554e-11 luc=-7.112508390e-18 wuc=2.584939414e-32 puc=-3.231174268e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.354238417e+05 lvsat=-1.382975091e-2 a0=-1.533380897e-02 la0=1.507103985e-7 ags=2.122259360e+00 lags=-1.472984367e-7 a1=0.0 a2=9.101975611e-01 la2=-2.727313031e-8 b0=0.0 b1=0.0 keta=-7.777436513e-02 lketa=1.101342597e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.768355118e-01 lpclm=-9.467448044e-9 pdiblc1=5.241829513e-01 lpdiblc1=-2.855766128e-8 pdiblc2=2.628226065e-02 lpdiblc2=-4.229372224e-9 pdiblcb=1.765059758e+00 lpdiblcb=-4.904191263e-07 ppdiblcb=8.881784197e-28 drout=-6.083418313e-01 ldrout=2.716006894e-7 pscbe1=7.999088729e+08 lpscbe1=1.538864396e-2 pscbe2=1.774695567e-08 lpscbe2=-2.126477355e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025125765e+01 lbeta0=-3.203990428e-7 agidl=-2.497675849e-09 lagidl=5.966198302e-16 bgidl=1.818113540e+09 lbgidl=-1.381548262e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.157772404e+00 lkt1=-3.251427011e-07 pkt1=8.881784197e-28 kt2=-5.770354749e-02 lkt2=1.168160598e-9 at=1.875627065e+05 lat=-2.858676971e-02 wat=1.862645149e-15 ute=-1.682167421e+00 lute=2.024611778e-7 ua1=1.624877580e-10 lua1=3.166184703e-17 ub1=-3.030938486e-19 lub1=3.195421259e-26 uc1=-2.633424711e-10 luc1=3.952258331e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.161 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.3e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='1.343870657e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.551556026e-07 wvth0=-1.678940596e-06 pvth0=3.120646887e-13 k1=3.437067510e-01 lk1=1.353118157e-07 wk1=4.991269153e-07 pk1=-9.277271974e-14 k2=-2.895249654e+00 lk2=4.990948174e-07 wk2=1.841020019e-06 pk2=-3.421903909e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.620398257e+00 ldsub=9.394577079e-07 wdsub=3.465394364e-06 pdsub=-6.441128505e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.199033583e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.888986352e-06 wvoff=2.172280948e-05 pvoff=-4.037618599e-12 nfactor='-4.916688436e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.173376928e-05 wnfactor=3.383799988e-04 pnfactor=-6.289469037e-11 eta0=-9.990807933e+00 leta0=1.948067771e-06 weta0=7.185872498e-06 peta0=-1.335638121e-12 etab=-5.875667322e-01 letab=1.090527184e-07 wetab=4.022646806e-07 petab=-7.476893618e-14 u0=-3.426538519e-02 lu0=7.088167780e-09 wu0=2.614624186e-08 pu0=-4.859801974e-15 ua=-5.419001772e-09 lua=6.304070318e-16 wua=2.325393564e-15 pua=-4.322209017e-22 ub=5.923011869e-18 lub=-7.172651474e-25 wub=-2.645788761e-24 pub=4.917727569e-31 uc=4.392686841e-10 luc=-8.412496379e-17 wuc=-3.103132565e-16 puc=5.767792498e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.045871875e+06 lvsat=-1.844469561e-01 wvsat=-6.803727952e-01 pvsat=1.264608914e-7 a0=5.555902870e+00 la0=-8.696434747e-07 wa0=-3.207868729e-06 pa0=5.962465607e-13 ags=1.250000057e+00 lags=-8.980734378e-15 wags=-2.601666438e-15 pags=4.835811751e-22 a1=0.0 a2=7.800522124e+00 la2=-1.310723320e-06 wa2=-4.834888570e-06 pa2=8.986607385e-13 b0=0.0 b1=0.0 keta=1.830144399e+00 lketa=-3.425027225e-07 wketa=-1.263395917e-06 pketa=2.348273991e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.592526162e-01 lpclm=-7.152395213e-09 wpclm=-2.638315620e-08 ppclm=4.903837243e-15 pdiblc1=-5.851099153e+00 lpdiblc1=1.153541148e-06 wpdiblc1=4.255088126e-06 ppdiblc1=-7.908932300e-13 pdiblc2=3.108731910e-02 lpdiblc2=-5.548255762e-09 wpdiblc2=-2.046595435e-08 ppdiblc2=3.804006935e-15 pdiblcb=3.493143043e+01 lpdiblcb=-6.704422521e-06 wpdiblcb=-2.473072352e-05 ppdiblcb=4.596699581e-12 drout=1.000000036e+00 ldrout=-1.875079647e-15 wdrout=8.533254459e-14 pdrout=-1.586076337e-20 pscbe1=1.476796236e+08 lpscbe1=1.212467884e+02 wpscbe1=4.472452013e+02 ppscbe1=-8.312946557e-5 pscbe2=1.417570559e-07 lpscbe2=-2.539030536e-14 wpscbe2=-9.365767662e-14 ppscbe2=1.740815235e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-3.902194178e+00 lbeta0=2.278048748e-06 wbeta0=8.403078730e-06 pbeta0=-1.561880244e-12 agidl=-3.623997061e-07 lagidl=6.755167141e-14 wagidl=2.491790599e-13 pagidl=-4.631491186e-20 bgidl=1.000000367e+09 lbgidl=-6.008681488e-05 wbgidl=-6.621429443e-05 pbgidl=1.230725861e-11 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-2.203433340e+01 lkt1=3.952842164e-06 wkt1=1.458091979e-05 pkt1=-2.710155562e-12 kt2=-1.487385738e+00 lkt2=2.670207870e-07 wkt2=9.849642433e-07 pkt2=-1.830753039e-13 at=1.288639548e+06 lat=-2.361217281e-01 wat=-8.709864303e-01 pat=1.618902478e-7 ute=1.036607634e+01 lute=-2.016564294e-06 wute=-7.438536998e-06 pute=1.382600872e-12 ua1=1.369256582e-08 lua1=-2.479986390e-15 wua1=-9.147969564e-15 pua1=1.700333103e-21 ub1=-1.819992810e-17 lub1=3.361655598e-24 wub1=1.240019885e-23 pub1=-2.304824961e-30 uc1=-4.392397940e-10 luc1=7.619532374e-17 wuc1=2.810630581e-16 puc1=-5.224119061e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.162 pmos lmin=2.0e-05 lmax=0.0001 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.163 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108621813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.532455644e-7 k1=4.171052081e-01 lk1=2.908460917e-7 k2=2.159455618e-02 lk2=-4.690448662e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=2.117582368e-27 pcit=4.743384505e-32 voff='-1.195937276e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.467000666e-6 nfactor='1.337826924e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.841077327e-5 eta0=0.08 etab=-0.07 u0=1.149534990e-02 lu0=-1.176644632e-8 ua=-9.044296180e-10 lua=2.075453526e-15 ub=1.700362603e-18 lub=-5.753769297e-24 wub=1.540743956e-39 uc=-1.046578370e-10 luc=-2.009187197e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.286628951e+04 lvsat=-2.540643246e-1 a0=1.625827411e+00 la0=-3.234747073e-6 ags=1.127460711e-01 lags=1.087252350e-8 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=-2.220025651e-07 lb0=2.392719013e-12 wb0=-1.058791184e-28 pb0=-8.470329473e-34 b1=-1.256728575e-09 lb1=2.383741859e-14 wb1=-3.101927297e-31 pb1=-6.617444900e-36 keta=3.416681995e-02 lketa=-2.159909532e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 wpclm=-2.775557562e-23 ppclm=6.661338148e-28 pdiblc1=0.39 pdiblc2=1.906905271e-03 lpdiblc2=-1.258792035e-8 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=8.865952071e-09 lpscbe2=2.388016187e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.797495750e+01 lbeta0=-3.592990887e-4 agidl=2.567367474e-09 lagidl=-1.413111313e-14 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.443649873e-01 lkt1=1.222316870e-07 wkt1=-4.440892099e-22 kt2=-6.519461656e-02 lkt2=1.328983321e-7 at=7.713361212e+04 lat=-1.228038641e-1 ute=5.595779957e-01 lute=-1.284400824e-05 wute=-2.220446049e-22 pute=4.440892099e-27 ua1=3.768264800e-09 lua1=-3.354261913e-14 ub1=-2.642787222e-18 lub1=2.826200788e-23 pub1=1.232595164e-44 uc1=-9.417115820e-11 luc1=1.286926591e-15 wuc1=-5.169878828e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.164 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.068786972e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.501020040e-8 k1=4.603509166e-01 lk1=-5.463825109e-8 k2=1.538364979e-02 lk2=2.713637080e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.472873697e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.816818865e-7 nfactor='9.225338883e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.233552538e-6 eta0=0.08 etab=-0.07 u0=8.814647214e-03 lu0=9.649338941e-9 ua=-8.481377777e-10 lua=1.625745332e-15 ub=1.054996270e-18 lub=-5.980215607e-25 uc=-1.070085284e-10 luc=-1.312504100e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.342054363e+04 lvsat=-1.882608877e-2 a0=1.169648264e+00 la0=4.096088288e-7 ags=4.536500838e-02 lags=5.491710742e-7 a1=0.0 a2=0.8 b0=5.791366221e-08 lb0=1.565046618e-13 b1=-1.307449963e-08 lb1=1.182480552e-13 pb1=2.646977960e-35 keta=7.536869066e-03 lketa=-3.247737421e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.061808156e-01 lpclm=4.371028699e-06 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=2.327209668e-04 lpdiblc2=7.869204170e-10 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.461096001e-08 lpscbe2=-2.201595970e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.997217500e-10 lalpha0=-7.966640969e-16 alpha1=1.997217500e-10 lalpha1=-7.966640969e-16 beta0=-2.392487250e+01 lbeta0=2.150993062e-4 agidl=4.330612791e-10 lagidl=2.919581601e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.139217330e-01 lkt1=-1.209755144e-7 kt2=-3.860015032e-02 lkt2=-7.956140140e-8 at=2.264263863e+04 lat=3.125174394e-1 ute=-1.910932237e+00 lute=6.892576840e-06 pute=7.105427358e-27 ua1=-2.943994399e-09 lua1=2.008074701e-14 ub1=2.913039917e-18 lub1=-1.612277288e-23 uc1=5.506278879e-10 luc1=-3.864289165e-15 wuc1=-1.033975766e-31 puc1=-1.654361225e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.165 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.063485550e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.386351842e-8 k1=3.863911154e-01 lk1=2.403777808e-7 k2=3.756574616e-02 lk2=-8.576786165e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.583304901e-01 ldsub=-1.190001542e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.285878909e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.082050964e-7 nfactor='8.585504846e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.681337744e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391132325e-01 letab=2.756836997e-7 u0=1.129776754e-02 lu0=-2.555052396e-10 ua=-3.948101738e-10 lua=-1.825195469e-16 ub=9.047694627e-19 lub=1.213642946e-27 uc=-1.333555795e-10 luc=1.037824576e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.345823238e+04 lvsat=-9.875382428e-2 a0=1.398566000e+00 la0=-5.035142625e-7 ags=-4.042771799e-02 lags=8.913871067e-7 a1=0.0 a2=0.8 b0=7.857195976e-08 lb0=7.410139848e-14 b1=2.737045909e-08 lb1=-4.308162726e-14 keta=2.253544784e-02 lketa=-6.307511832e-08 wketa=-1.387778781e-23 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.074223900e-01 lpclm=3.278972801e-7 pdiblc1=0.39 pdiblc2=4.187393462e-04 lpdiblc2=4.491728403e-11 pdiblcb=-4.238870000e-01 lpdiblcb=7.933343877e-7 drout=0.56 pscbe1=800000000.0 pscbe2=8.718970657e-09 lpscbe2=1.486419869e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-9.944350000e-11 lalpha0=3.966671938e-16 alpha1=-9.944350000e-11 lalpha1=3.966671938e-16 beta0=5.429614004e+01 lbeta0=-9.691414411e-5 agidl=9.014407177e-10 lagidl=1.051276909e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.356779703e-01 lkt1=-3.419271211e-8 kt2=-6.313133978e-02 lkt2=1.829032431e-8 at=1.615988244e+05 lat=-2.417607213e-1 ute=-9.311290905e-02 lute=-3.584681431e-7 ua1=2.873317563e-09 lua1=-3.123754152e-15 ub1=-1.891532202e-18 lub1=3.042040710e-24 uc1=-8.692813487e-10 luc1=1.799544192e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.166 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.081024143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.874549914e-8 k1=5.064919019e-01 lk1=1.512929702e-9 k2=-5.250837621e-03 lk2=-6.112426770e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.600000199e-01 ldsub=-1.966733887e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.854733267e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.224558331e-7 nfactor='7.974519768e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.466167851e-6 eta0=-4.835518650e-01 leta0=9.627162327e-07 weta0=-3.122502257e-23 peta0=3.747002708e-28 etab=2.386594872e-04 letab=-1.469097694e-9 u0=1.277578903e-02 lu0=-3.195097838e-9 ua=-2.787126111e-10 lua=-4.134225064e-16 ub=8.338866336e-19 lub=1.421903751e-25 uc=-1.183445084e-10 luc=7.392738859e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.599790864e+04 lvsat=3.541598979e-2 a0=1.034813481e+00 la0=2.199422095e-7 ags=2.529917783e-01 lags=3.078138731e-7 a1=0.0 a2=0.8 b0=1.262823559e-07 lb0=-2.078837708e-14 b1=9.908435342e-09 lb1=-8.351932082e-15 keta=-1.722971284e-02 lketa=1.601261680e-08 wketa=-1.387778781e-23 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.149196182e-01 lpclm=-2.836747322e-07 wpclm=-8.881784197e-22 pdiblc1=3.955978546e-01 lpdiblc1=-1.113340513e-8 pdiblc2=4.525213076e-04 lpdiblc2=-2.227064540e-11 pdiblcb=1.727740000e-01 lpdiblcb=-3.933467754e-07 ppdiblcb=-1.110223025e-28 drout=3.855974777e-01 ldrout=3.468639446e-7 pscbe1=800000000.0 pscbe2=9.759262277e-09 lpscbe2=-5.825849256e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.674544110e+00 lbeta0=1.776759381e-6 agidl=1.018141354e-09 lagidl=8.191745147e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.269668075e-01 lkt1=-5.151808255e-8 kt2=-5.925098613e-02 lkt2=1.057280534e-8 at=2.845269774e+04 lat=2.304961559e-2 ute=4.928361669e-01 lute=-1.523844682e-6 ua1=3.016514543e-09 lua1=-3.408554329e-15 ub1=-1.565341614e-18 lub1=2.393290035e-24 uc1=4.482619664e-12 luc1=6.174124785e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.167 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.054442900e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.246010562e-8 k1=5.794701714e-01 lk1=-7.065309168e-8 k2=-3.599095491e-02 lk2=2.978673710e-08 wk2=-6.938893904e-24 pk2=1.040834086e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.635276000e-01 ldsub=7.154747378e-07 pdsub=-2.220446049e-28 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.984410505e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.639222613e-8 nfactor='8.580472176e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.065376009e-6 eta0=9.611039418e-01 leta0=-4.658605549e-7 etab=-1.488450021e-03 letab=2.387890846e-10 u0=-3.953040131e-03 lu0=1.334753945e-08 pu0=6.938893904e-30 ua=-2.555715282e-09 lua=1.838237125e-15 wua=-8.271806126e-31 pua=8.271806126e-37 ub=1.635833473e-19 lub=8.050331859e-25 uc=-3.894326448e-11 luc=-4.590119479e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.069252850e+04 lvsat=1.107521054e-3 a0=1.396980751e+00 la0=-1.381941390e-7 ags=-1.061952942e-01 lags=6.630031935e-7 a1=0.0 a2=1.100991363e+00 la2=-2.976413294e-07 wa2=-8.881784197e-22 b0=2.081769124e-07 lb0=-1.017714472e-13 b1=2.892444750e-09 lb1=-1.414029465e-15 keta=4.051134126e-02 lketa=-4.108577937e-08 wketa=1.734723476e-24 pketa=8.673617380e-30 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=8.192448538e-01 lpclm=-1.890648279e-7 pdiblc1=6.918059423e-01 lpdiblc1=-3.040446968e-07 wpdiblc1=-4.440892099e-22 pdiblc2=6.468668115e-05 lpdiblc2=3.612473816e-10 pdiblcb=-0.225 drout=9.557609593e-01 ldrout=-2.169536175e-07 wdrout=-8.881784197e-22 pscbe1=1.446985488e+09 lpscbe1=-6.397845396e+02 ppscbe1=4.768371582e-19 pscbe2=-5.829857018e-08 lpscbe2=6.671776386e-14 ppscbe2=-2.646977960e-35 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.544352635e+00 lbeta0=1.905501825e-6 agidl=1.849125933e-09 lagidl=-2.561206190e-18 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.743566677e-01 lkt1=-4.655671468e-9 kt2=-3.781888407e-02 lkt2=-1.062075742e-8 at=2.415206960e+04 lat=2.730237773e-2 ute=-1.839698799e+00 lute=7.827291698e-7 ua1=-2.479750931e-09 lua1=2.026537710e-15 pua1=-4.135903063e-37 ub1=2.537894393e-18 lub1=-1.664276955e-24 uc1=1.981977632e-10 luc1=-1.298178461e-16 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.168 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.795119211e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.417140212e-8 k1=2.983925622e-01 lk1=6.675731910e-8 k2=6.116802299e-02 lk2=-1.771137242e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.205819134e+00 ldsub=-1.006188000e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.202390991e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.704863814e-8 nfactor='4.297447230e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.846639641e-8 eta0=-4.522078841e-01 leta0=2.250651974e-07 weta0=-1.526556659e-22 peta0=-5.204170428e-29 etab=-1.886870119e-03 letab=4.335647182e-10 u0=3.805558220e-02 lu0=-7.189215745e-9 ua=3.372214182e-09 lua=-1.059749752e-15 pua=-4.135903063e-37 ub=1.910230175e-18 lub=-4.885004854e-26 uc=-9.356751888e-11 luc=2.211403977e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.948254123e+04 lvsat=1.147644753e-2 a0=1.590800918e+00 la0=-2.329470036e-7 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=2.018182291e-01 la2=1.419374407e-7 b0=0.0 b1=0.0 keta=-5.486585336e-02 lketa=5.541269763e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.369246124e-01 lpclm=9.561406851e-8 pdiblc1=-2.499817842e-01 lpdiblc1=1.563670691e-07 wpdiblc1=-1.110223025e-22 ppdiblc1=5.551115123e-29 pdiblc2=-6.623202468e-03 lpdiblc2=3.630755750e-09 wpdiblc2=-1.734723476e-24 ppdiblc2=-6.505213035e-31 pdiblcb=-1.647857919e-01 lpdiblcb=-2.943691991e-8 drout=4.960126660e-01 ldrout=7.803530650e-9 pscbe1=-4.939454606e+08 lpscbe1=3.090783733e+02 ppscbe1=5.960464478e-20 pscbe2=1.444184156e-07 lpscbe2=-3.238448899e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=7.995122502e+00 lbeta0=2.185239603e-7 agidl=3.605683955e-09 lagidl=-8.612897264e-16 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.518752346e-01 lkt1=1.310148304e-7 kt2=-6.597515796e-02 lkt2=3.144000191e-9 at=9.157306403e+04 lat=-5.657723812e-3 ute=3.308550878e-01 lute=-2.783895088e-07 pute=1.110223025e-28 ua1=2.975146297e-09 lua1=-6.401978981e-16 ub1=-1.532522831e-18 lub1=3.256279136e-25 uc1=-3.817149149e-11 luc1=-1.426400859e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.169 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.794369863e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.807630180e-8 k1=-6.134766510e-01 lk1=2.845755181e-7 k2=4.624846070e-01 lk2=-1.135738648e-07 wk2=5.551115123e-23 pk2=-2.775557562e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.630409017e+00 ldsub=-2.020405853e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.038439192e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.701932152e-8 nfactor='1.056398954e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.468422564e-6 eta0=4.900000007e-01 leta0=-5.142020143e-17 etab=1.809698392e-03 letab=-4.494346021e-10 wetab=8.673617380e-25 petab=1.355252716e-31 u0=1.782350564e-02 lu0=-2.356379616e-9 ua=1.258985607e-09 lua=-5.549628425e-16 ub=8.412917613e-19 lub=2.064872702e-25 uc=2.878584554e-11 luc=-7.112508390e-18 wuc=9.693522803e-33 puc=-1.615587134e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.354238417e+05 lvsat=-1.382975091e-2 a0=-1.533380897e-02 la0=1.507103985e-7 ags=2.122259360e+00 lags=-1.472984367e-7 a1=0.0 a2=9.101975611e-01 la2=-2.727313031e-8 b0=0.0 b1=0.0 keta=-7.777436513e-02 lketa=1.101342597e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.768355118e-01 lpclm=-9.467448044e-9 pdiblc1=5.241829513e-01 lpdiblc1=-2.855766128e-8 pdiblc2=2.628226065e-02 lpdiblc2=-4.229372224e-9 pdiblcb=1.765059758e+00 lpdiblcb=-4.904191263e-07 wpdiblcb=-8.881784197e-22 drout=-6.083418313e-01 ldrout=2.716006894e-7 pscbe1=7.999088729e+08 lpscbe1=1.538864396e-2 pscbe2=1.774695567e-08 lpscbe2=-2.126477355e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025125765e+01 lbeta0=-3.203990428e-7 agidl=-2.497675849e-09 lagidl=5.966198302e-16 bgidl=1.818113540e+09 lbgidl=-1.381548262e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.157772404e+00 lkt1=-3.251427011e-07 pkt1=-1.110223025e-28 kt2=-5.770354749e-02 lkt2=1.168160598e-9 at=1.875627065e+05 lat=-2.858676971e-02 pat=2.910383046e-23 ute=-1.682167421e+00 lute=2.024611778e-7 ua1=1.624877580e-10 lua1=3.166184703e-17 ub1=-3.030938486e-19 lub1=3.195421259e-26 uc1=-2.633424711e-10 luc1=3.952258331e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.170 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=6.3e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.093926099e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.042319483e-09 wvth0=-3.191147638e-08 pvth0=5.931386115e-15 k1=3.319605812e-01 lk1=1.374950763e-07 wk1=5.070628860e-07 pk1=-9.424777862e-14 k2=3.144826514e-01 lk2=-9.749812623e-08 wk2=-3.275457409e-07 pk2=6.088092686e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.701950988e+00 ldsub=9.546159140e-07 wdsub=3.520493183e-06 pdsub=-6.543540680e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='4.563649242e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-9.053028539e-07 wvoff=-2.973867019e-06 pvoff=5.527526629e-13 nfactor='6.259221849e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.128673434e-05 wnfactor=-3.609096854e-05 pnfactor=6.708228323e-12 eta0=-9.990807256e+00 leta0=1.948067645e-06 weta0=7.185872041e-06 peta0=-1.335638036e-12 etab=-5.970333503e-01 letab=1.108122787e-07 wetab=4.086605360e-07 petab=-7.595773382e-14 u0=2.161004568e-03 lu0=3.175947159e-10 wu0=1.535771558e-09 pu0=-2.854538595e-16 ua=-5.418884288e-09 lua=6.303851951e-16 wua=2.325314189e-15 pua=-4.322061483e-22 ub=5.923003290e-18 lub=-7.172635528e-25 wub=-2.645782964e-24 pub=4.917716796e-31 uc=4.465714238e-10 luc=-8.548232402e-17 wuc=-3.152471481e-16 puc=5.859498742e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.914692273e+05 lvsat=8.271163450e-02 wvsat=2.907264748e-01 pvsat=-5.403732987e-8 a0=5.555903394e+00 la0=-8.696435721e-07 wa0=-3.207869083e-06 pa0=5.962466265e-13 ags=1.250000053e+00 lags=-8.187253542e-15 wags=2.825188972e-16 pags=-5.251177271e-23 a1=0.0 a2=7.914304040e+00 la2=-1.331871965e-06 wa2=-4.911762136e-06 pa2=9.129492282e-13 b0=0.0 b1=0.0 keta=1.830144754e+00 lketa=-3.425027884e-07 wketa=-1.263396156e-06 pketa=2.348274436e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.598735084e-01 lpclm=-7.267800440e-09 wpclm=-2.680264461e-08 ppclm=4.981807553e-15 pdiblc1=-5.951236129e+00 lpdiblc1=1.172153608e-06 wpdiblc1=4.322742870e-06 ppdiblc1=-8.034682172e-13 pdiblc2=3.156894820e-02 lpdiblc2=-5.637776163e-09 wpdiblc2=-2.079135357e-08 ppdiblc2=3.864488888e-15 pdiblcb=3.551343339e+01 lpdiblcb=-6.812599412e-06 wpdiblcb=-2.512393753e-05 ppdiblcb=4.669786268e-12 drout=1.000000176e+00 ldrout=-2.790014442e-14 wdrout=-9.266393874e-15 pdrout=1.722344045e-21 pscbe1=1.371544465e+08 lpscbe1=1.232031030e+02 wpscbe1=4.543562426e+02 ppscbe1=-8.445119480e-5 pscbe2=1.439611197e-07 lpscbe2=-2.579997469e-14 wpscbe2=-9.514679060e-14 ppscbe2=1.768493397e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-4.099948165e+00 lbeta0=2.314805282e-06 wbeta0=8.536685675e-06 pbeta0=-1.586713766e-12 agidl=4.780010855e-08 lagidl=-8.692168143e-15 wagidl=-2.796095931e-14 pagidl=5.197103506e-21 bgidl=1.000000258e+09 lbgidl=-3.989249611e-05 wbgidl=7.190319061e-06 pbgidl=-1.336463928e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.184876322e-01 lkt1=-8.348208875e-08 wkt1=-9.078335883e-08 pkt1=1.687390291e-14 kt2=-1.510565206e+00 lkt2=2.713291548e-07 wkt2=1.000624802e-06 pkt2=-1.859861320e-13 at=1.309136784e+06 lat=-2.399315494e-01 wat=-8.848348139e-01 pat=1.644642469e-7 ute=1.054113156e+01 lute=-2.049101809e-06 wute=-7.556808160e-06 pute=1.404583933e-12 ua1=1.390785269e-08 lua1=-2.520001761e-15 wua1=-9.293422110e-15 pua1=1.727368368e-21 ub1=-1.849174368e-17 lub1=3.415895360e-24 wub1=1.259735588e-23 pub1=-2.341470537e-30 uc1=-4.458541873e-10 luc1=7.742474102e-17 wuc1=2.855318877e-16 puc1=-5.307181197e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.171 pmos lmin=2.0e-05 lmax=0.0001 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.172 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.108621813e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.532455644e-07 wvth0=7.105427358e-21 k1=4.171052081e-01 lk1=2.908460917e-7 k2=2.159455618e-02 lk2=-4.690448662e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=1.355252716e-26 pcit=1.084202172e-31 voff='-1.195937276e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.467000666e-6 nfactor='1.337826924e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.841077327e-5 eta0=0.08 etab=-0.07 u0=1.149534990e-02 lu0=-1.176644632e-8 ua=-9.044296180e-10 lua=2.075453526e-15 ub=1.700362603e-18 lub=-5.753769297e-24 uc=-1.046578370e-10 luc=-2.009187197e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.286628951e+04 lvsat=-2.540643246e-1 a0=1.625827411e+00 la0=-3.234747073e-6 ags=1.127460711e-01 lags=1.087252350e-8 a1=0.0 a2=1.083175658e+00 la2=-2.262253522e-6 b0=-2.220025651e-07 lb0=2.392719013e-12 wb0=-8.470329473e-28 b1=-1.256728575e-09 lb1=2.383741859e-14 wb1=-2.481541838e-30 pb1=-4.632211430e-35 keta=3.416681995e-02 lketa=-2.159909532e-7 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-6.885582638e-02 lpclm=1.676183212e-06 wpclm=-1.110223025e-22 ppclm=3.552713679e-27 pdiblc1=0.39 pdiblc2=1.906905271e-03 lpdiblc2=-1.258792035e-8 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=8.865952071e-09 lpscbe2=2.388016187e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-6.657391667e-11 lalpha0=1.330737366e-15 alpha1=-6.657391667e-11 lalpha1=1.330737366e-15 beta0=4.797495750e+01 lbeta0=-3.592990887e-4 agidl=2.567367474e-09 lagidl=-1.413111313e-14 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.443649873e-01 lkt1=1.222316870e-7 kt2=-6.519461656e-02 lkt2=1.328983321e-7 at=7.713361212e+04 lat=-1.228038641e-1 ute=5.595779957e-01 lute=-1.284400824e-05 pute=-1.421085472e-26 ua1=3.768264800e-09 lua1=-3.354261913e-14 ub1=-2.642787222e-18 lub1=2.826200788e-23 pub1=9.860761315e-44 uc1=-9.417115820e-11 luc1=1.286926591e-15 puc1=3.308722450e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.173 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.068786972e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.501020040e-8 k1=4.603509166e-01 lk1=-5.463825109e-8 k2=1.538364979e-02 lk2=2.713637080e-9 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.472873697e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.816818865e-7 nfactor='9.225338883e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-5.233552538e-6 eta0=0.08 etab=-0.07 u0=8.814647214e-03 lu0=9.649338941e-9 ua=-8.481377777e-10 lua=1.625745332e-15 ub=1.054996270e-18 lub=-5.980215607e-25 uc=-1.070085284e-10 luc=-1.312504100e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.342054363e+04 lvsat=-1.882608877e-2 a0=1.169648264e+00 la0=4.096088288e-7 ags=4.536500838e-02 lags=5.491710742e-7 a1=0.0 a2=0.8 b0=5.791366221e-08 lb0=1.565046618e-13 b1=-1.307449963e-08 lb1=1.182480552e-13 pb1=-3.176373552e-34 keta=7.536869066e-03 lketa=-3.247737421e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.061808156e-01 lpclm=4.371028699e-6 pdiblc1=0.39 pdiblc2=2.327209668e-04 lpdiblc2=7.869204170e-10 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.461096001e-08 lpscbe2=-2.201595970e-14 wpscbe2=-1.058791184e-28 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.997217500e-10 lalpha0=-7.966640969e-16 alpha1=1.997217500e-10 lalpha1=-7.966640969e-16 beta0=-2.392487250e+01 lbeta0=2.150993062e-04 wbeta0=2.842170943e-20 pbeta0=-3.410605132e-25 agidl=4.330612791e-10 lagidl=2.919581601e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.139217330e-01 lkt1=-1.209755144e-7 kt2=-3.860015032e-02 lkt2=-7.956140140e-8 at=2.264263863e+04 lat=3.125174394e-1 ute=-1.910932237e+00 lute=6.892576840e-6 ua1=-2.943994399e-09 lua1=2.008074701e-14 wua1=-6.617444900e-30 pua1=2.646977960e-35 ub1=2.913039917e-18 lub1=-1.612277288e-23 uc1=5.506278879e-10 luc1=-3.864289165e-15 wuc1=-1.654361225e-30 puc1=9.926167351e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.174 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.063485550e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.386351842e-8 k1=3.863911154e-01 lk1=2.403777808e-7 k2=3.756574616e-02 lk2=-8.576786165e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.583304901e-01 ldsub=-1.190001542e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.285878909e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.082050964e-7 nfactor='8.585504846e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.681337744e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391132325e-01 letab=2.756836997e-7 u0=1.129776754e-02 lu0=-2.555052396e-10 ua=-3.948101738e-10 lua=-1.825195469e-16 ub=9.047694627e-19 lub=1.213642946e-27 uc=-1.333555795e-10 luc=1.037824576e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.345823238e+04 lvsat=-9.875382428e-2 a0=1.398566000e+00 la0=-5.035142625e-7 ags=-4.042771799e-02 lags=8.913871067e-7 a1=0.0 a2=0.8 b0=7.857195976e-08 lb0=7.410139848e-14 b1=2.737045909e-08 lb1=-4.308162726e-14 keta=2.253544784e-02 lketa=-6.307511832e-08 wketa=5.551115123e-23 pketa=1.110223025e-28 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.074223900e-01 lpclm=3.278972801e-7 pdiblc1=0.39 pdiblc2=4.187393462e-04 lpdiblc2=4.491728403e-11 pdiblcb=-4.238870000e-01 lpdiblcb=7.933343877e-7 drout=0.56 pscbe1=800000000.0 pscbe2=8.718970657e-09 lpscbe2=1.486419869e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-9.944350000e-11 lalpha0=3.966671938e-16 alpha1=-9.944350000e-11 lalpha1=3.966671938e-16 beta0=5.429614004e+01 lbeta0=-9.691414411e-5 agidl=9.014407177e-10 lagidl=1.051276909e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.356779703e-01 lkt1=-3.419271211e-8 kt2=-6.313133979e-02 lkt2=1.829032431e-8 at=1.615988244e+05 lat=-2.417607213e-1 ute=-9.311290905e-02 lute=-3.584681431e-7 ua1=2.873317562e-09 lua1=-3.123754152e-15 ub1=-1.891532202e-18 lub1=3.042040710e-24 uc1=-8.692813487e-10 luc1=1.799544192e-15 puc1=6.617444900e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.175 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.081024143e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=4.874549914e-8 k1=5.064919019e-01 lk1=1.512929702e-9 k2=-5.250837621e-03 lk2=-6.112426770e-10 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=2.600000199e-01 ldsub=-1.966733620e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.854733267e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=1.224558331e-7 nfactor='7.974519768e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.466167851e-6 eta0=-4.835518650e-01 leta0=9.627162327e-07 weta0=-8.118505868e-22 peta0=2.851885395e-27 etab=2.386594872e-04 letab=-1.469097694e-9 u0=1.277578903e-02 lu0=-3.195097838e-9 ua=-2.787126111e-10 lua=-4.134225064e-16 ub=8.338866336e-19 lub=1.421903751e-25 uc=-1.183445084e-10 luc=7.392738859e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.599790864e+04 lvsat=3.541598979e-2 a0=1.034813481e+00 la0=2.199422095e-7 ags=2.529917783e-01 lags=3.078138731e-7 a1=0.0 a2=0.8 b0=1.262823559e-07 lb0=-2.078837708e-14 b1=9.908435342e-09 lb1=-8.351932082e-15 keta=-1.722971284e-02 lketa=1.601261680e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.149196182e-01 lpclm=-2.836747322e-7 pdiblc1=3.955978546e-01 lpdiblc1=-1.113340513e-8 pdiblc2=4.525213076e-04 lpdiblc2=-2.227064540e-11 pdiblcb=1.727740000e-01 lpdiblcb=-3.933467754e-07 wpdiblcb=-2.220446049e-22 ppdiblcb=-4.440892099e-28 drout=3.855974777e-01 ldrout=3.468639446e-7 pscbe1=800000000.0 pscbe2=9.759262277e-09 lpscbe2=-5.825849256e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.674544110e+00 lbeta0=1.776759381e-6 agidl=1.018141354e-09 lagidl=8.191745147e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.269668075e-01 lkt1=-5.151808255e-8 kt2=-5.925098613e-02 lkt2=1.057280534e-8 at=2.845269774e+04 lat=2.304961559e-2 ute=4.928361669e-01 lute=-1.523844682e-6 ua1=3.016514543e-09 lua1=-3.408554329e-15 ub1=-1.565341614e-18 lub1=2.393290035e-24 wub1=-3.081487911e-39 uc1=4.482619664e-12 luc1=6.174124785e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.176 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.054442900e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.246010562e-8 k1=5.794701714e-01 lk1=-7.065309168e-8 k2=-3.599095491e-02 lk2=2.978673710e-08 wk2=-5.551115123e-23 pk2=8.326672685e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.635276000e-01 ldsub=7.154747378e-07 pdsub=-1.776356839e-27 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.984410505e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.639222613e-8 nfactor='8.580472176e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.065376009e-6 eta0=9.611039418e-01 leta0=-4.658605549e-7 etab=-1.488450021e-03 letab=2.387890846e-10 u0=-3.953040131e-03 lu0=1.334753945e-8 ua=-2.555715282e-09 lua=1.838237125e-15 wua=6.617444900e-30 pua=3.308722450e-36 ub=1.635833473e-19 lub=8.050331859e-25 uc=-3.894326448e-11 luc=-4.590119479e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.069252850e+04 lvsat=1.107521054e-3 a0=1.396980751e+00 la0=-1.381941390e-7 ags=-1.061952942e-01 lags=6.630031935e-7 a1=0.0 a2=1.100991363e+00 la2=-2.976413294e-7 b0=2.081769124e-07 lb0=-1.017714472e-13 b1=2.892444750e-09 lb1=-1.414029465e-15 keta=4.051134126e-02 lketa=-4.108577937e-08 wketa=9.714451465e-23 pketa=5.551115123e-29 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=8.192448538e-01 lpclm=-1.890648279e-7 pdiblc1=6.918059423e-01 lpdiblc1=-3.040446968e-7 pdiblc2=6.468668115e-05 lpdiblc2=3.612473816e-10 pdiblcb=-0.225 drout=9.557609593e-01 ldrout=-2.169536175e-7 pscbe1=1.446985488e+09 lpscbe1=-6.397845396e+2 pscbe2=-5.829857018e-08 lpscbe2=6.671776386e-14 wpscbe2=-1.058791184e-28 ppscbe2=-2.117582368e-34 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=4.544352635e+00 lbeta0=1.905501825e-6 agidl=1.849125933e-09 lagidl=-2.561206190e-18 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.743566677e-01 lkt1=-4.655671468e-9 kt2=-3.781888407e-02 lkt2=-1.062075742e-8 at=2.415206960e+04 lat=2.730237773e-2 ute=-1.839698799e+00 lute=7.827291698e-7 ua1=-2.479750931e-09 lua1=2.026537710e-15 pua1=-1.654361225e-36 ub1=2.537894393e-18 lub1=-1.664276955e-24 uc1=1.981977632e-10 luc1=-1.298178461e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.177 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.795119211e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.417140212e-8 k1=2.983925622e-01 lk1=6.675731910e-8 k2=6.116802299e-02 lk2=-1.771137242e-08 wk2=2.220446049e-22 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.205819134e+00 ldsub=-1.006188000e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.202390991e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.704863814e-8 nfactor='4.297447230e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.846639641e-8 eta0=-4.522078841e-01 leta0=2.250651974e-07 weta0=-7.771561172e-22 peta0=8.326672685e-29 etab=-1.886870119e-03 letab=4.335647182e-10 u0=3.805558220e-02 lu0=-7.189215745e-9 ua=3.372214182e-09 lua=-1.059749752e-15 wua=-1.323488980e-29 ub=1.910230175e-18 lub=-4.885004854e-26 uc=-9.356751888e-11 luc=2.211403977e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.948254123e+04 lvsat=1.147644753e-2 a0=1.590800918e+00 la0=-2.329470036e-7 ags=1.005767373e+00 lags=1.193980042e-7 a1=0.0 a2=2.018182291e-01 la2=1.419374407e-7 b0=0.0 b1=0.0 keta=-5.486585336e-02 lketa=5.541269763e-9 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.369246124e-01 lpclm=9.561406851e-8 pdiblc1=-2.499817842e-01 lpdiblc1=1.563670691e-07 wpdiblc1=8.881784197e-22 ppdiblc1=-2.220446049e-28 pdiblc2=-6.623202468e-03 lpdiblc2=3.630755750e-09 wpdiblc2=-6.938893904e-24 ppdiblc2=-1.040834086e-29 pdiblcb=-1.647857919e-01 lpdiblcb=-2.943691991e-8 drout=4.960126660e-01 ldrout=7.803530650e-9 pscbe1=-4.939454606e+08 lpscbe1=3.090783733e+02 wpscbe1=-1.907348633e-12 ppscbe1=9.536743164e-19 pscbe2=1.444184156e-07 lpscbe2=-3.238448899e-14 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=7.995122502e+00 lbeta0=2.185239603e-7 agidl=3.605683955e-09 lagidl=-8.612897264e-16 bgidl=7.709281792e+08 lbgidl=1.119863410e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=-7.518752346e-01 lkt1=1.310148304e-7 kt2=-6.597515796e-02 lkt2=3.144000191e-9 at=9.157306403e+04 lat=-5.657723812e-3 ute=3.308550878e-01 lute=-2.783895088e-07 pute=-4.440892099e-28 ua1=2.975146297e-09 lua1=-6.401978981e-16 ub1=-1.532522831e-18 lub1=3.256279136e-25 uc1=-3.817149149e-11 luc1=-1.426400859e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.178 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-8.794369863e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-3.807630180e-8 k1=-6.134766510e-01 lk1=2.845755181e-7 k2=4.624846070e-01 lk2=-1.135738648e-07 wk2=8.881784197e-22 pk2=5.551115123e-29 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.630409017e+00 ldsub=-2.020405853e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.038439192e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.701932152e-8 nfactor='1.056398954e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.468422564e-6 eta0=4.900000007e-01 leta0=-5.141842507e-17 etab=1.809698392e-03 letab=-4.494346021e-10 wetab=-5.204170428e-24 petab=-1.084202172e-30 u0=1.782350564e-02 lu0=-2.356379616e-9 ua=1.258985607e-09 lua=-5.549628425e-16 ub=8.412917613e-19 lub=2.064872702e-25 uc=2.878584554e-11 luc=-7.112508390e-18 wuc=-5.169878828e-32 puc=-1.615587134e-38 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.354238417e+05 lvsat=-1.382975091e-2 a0=-1.533380897e-02 la0=1.507103985e-7 ags=2.122259360e+00 lags=-1.472984367e-7 a1=0.0 a2=9.101975611e-01 la2=-2.727313031e-8 b0=0.0 b1=0.0 keta=-7.777436513e-02 lketa=1.101342597e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.768355118e-01 lpclm=-9.467448044e-9 pdiblc1=5.241829513e-01 lpdiblc1=-2.855766128e-8 pdiblc2=2.628226065e-02 lpdiblc2=-4.229372224e-9 pdiblcb=1.765059758e+00 lpdiblcb=-4.904191263e-07 ppdiblcb=8.881784197e-28 drout=-6.083418313e-01 ldrout=2.716006894e-7 pscbe1=7.999088729e+08 lpscbe1=1.538864396e-2 pscbe2=1.774695567e-08 lpscbe2=-2.126477355e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.025125765e+01 lbeta0=-3.203990428e-7 agidl=-2.497675849e-09 lagidl=5.966198302e-16 bgidl=1.818113540e+09 lbgidl=-1.381548262e+2 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644019647032 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.29936672419988e-10 mjswgs=0.70393 tnom=30.0 kt1=1.157772404e+00 lkt1=-3.251427011e-7 kt2=-5.770354749e-02 lkt2=1.168160598e-9 at=1.875627065e+05 lat=-2.858676971e-2 ute=-1.682167421e+00 lute=2.024611778e-7 ua1=1.624877580e-10 lua1=3.166184703e-17 ub1=-3.030938486e-19 lub1=3.195421259e-26 uc1=-2.633424711e-10 luc1=3.952258331e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.179 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='4.543996377e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.049962970e-06 wvth0=-3.389982137e-06 pvth0=6.300959799e-13 k1=-2.258766977e-01 lk1=2.411802913e-07 wk1=8.393230418e-07 pk1=-1.560049738e-13 k2=-3.242967156e+00 lk2=5.637250696e-07 wk2=1.791349629e-06 pk2=-3.329581555e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=4.848290830e+00 ldsub=-8.204875327e-07 wdsub=-2.167840949e-06 pdsub=4.029365972e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.253162774e+01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.989596279e-06 wvoff=1.912089605e-05 pvoff=-3.554000949e-12 nfactor='-4.442400929e+02+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=8.291818738e-05 wnfactor=2.657895064e-04 pnfactor=-4.940229556e-11 eta0=7.745943157e+00 leta0=-1.348662154e-06 weta0=-3.378526713e-06 peta0=6.279667602e-13 etab=4.049986945e-01 letab=-7.543541751e-08 wetab=-1.881717946e-07 petab=3.497549146e-14 u0=-2.800481726e-02 lu0=5.924516019e-09 wu0=1.950319869e-08 pu0=-3.625059540e-15 ua=8.933726323e-09 lua=-2.037334539e-15 wua=-6.223416448e-15 pua=1.156746415e-21 ub=-1.166844130e-18 lub=6.005263871e-25 wub=1.577086136e-24 pub=-2.931330000e-31 uc=-4.282788327e-10 luc=7.712609314e-17 wuc=2.058329114e-16 puc=-3.825816323e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.550727464e+06 lvsat=-6.500244645e-01 wvsat=-2.057332603e+00 pvsat=3.823964109e-7 a0=2.201214274e-02 la0=1.589407948e-07 wa0=8.823829167e-08 pa0=-1.640085127e-14 ags=1.249999926e+00 lags=1.538647609e-14 wags=7.582468697e-14 pags=-1.409353700e-20 a1=0.0 a2=-6.144436002e+00 la2=1.281226047e-06 wa2=3.461932726e-06 pa2=-6.434694357e-13 b0=0.0 b1=0.0 keta=-1.375383862e+00 lketa=2.533088155e-07 wketa=6.458872091e-07 pketa=-1.200510555e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=6.628759095e-01 lpclm=-7.825856746e-09 wpclm=-2.859094080e-08 ppclm=5.314198166e-15 pdiblc1=1.148677440e+00 lpdiblc1=-1.475073275e-07 wpdiblc1=9.387815034e-08 ppdiblc1=-1.744913180e-14 pdiblc2=2.527577101e-02 lpdiblc2=-4.468063319e-09 wpdiblc2=-1.704299878e-08 ppdiblc2=3.167782184e-15 pdiblcb=-1.443754083e+01 lpdiblcb=2.471788166e-06 wpdiblcb=4.627961642e-06 ppdiblcb=-8.601992303e-13 drout=1.000000030e+00 ldrout=-8.456240153e-16 wdrout=7.743003039e-14 pdrout=-1.439192232e-20 pscbe1=1.246682778e+09 lpscbe1=-8.302492798e+01 wpscbe1=-2.065032415e+02 ppscbe1=3.838275749e-5 pscbe2=-1.060382373e-08 lpscbe2=2.929011338e-15 wpscbe2=-3.084509878e-15 ppscbe2=5.733178510e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.725114145e+01 lbeta0=-1.653721745e-06 wbeta0=-4.180493024e-06 pbeta0=7.770282384e-13 agidl=-3.246694584e-07 lagidl=6.053875026e-14 wagidl=1.938901091e-13 pagidl=-3.603835458e-20 bgidl=1.000000359e+09 lbgidl=-5.860388184e-05 wbgidl=-5.277047729e-05 pbgidl=9.808448792e-12 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=5.202529742e+00 lkt1=-1.109673588e-06 wkt1=-3.379222769e-06 pkt1=6.280961361e-13 kt2=9.691529664e-01 lkt2=-1.895760619e-07 wkt2=-4.763498952e-07 pkt2=8.853915502e-14 at=-5.116395771e+05 lat=9.849615283e-02 wat=1.996596437e-01 pat=-3.711073798e-8 ute=-2.146123259e+00 lute=3.090782449e-07 wute=-6.872357972e-14 pute=1.277365058e-20 ua1=1.104806946e-10 lua1=4.451577126e-17 wua1=-1.075403810e-15 pua1=1.998853061e-22 ub1=2.980863316e-18 lub1=-5.752181021e-25 wub1=-1.922012433e-25 pub1=3.572444508e-32 uc1=-7.122960440e-10 luc1=1.269482889e-16 wuc1=4.442305192e-16 puc1=-8.256912661e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.180 pmos lmin=2.0e-05 lmax=0.0001 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.181 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.142544781e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.031327361e-06 wvth0=1.986603635e-08 pvth0=-3.970996179e-13 k1=3.602134186e-01 lk1=1.428048676e-06 wk1=3.331708355e-08 pk1=-6.659708518e-13 k2=2.591525663e-02 lk2=-1.332704063e-07 wk2=-2.530297242e-09 pk2=5.057778264e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=6.352747104e-28 pcit=-1.863472484e-32 voff='-1.201320773e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.574610691e-06 wvoff=3.152694373e-09 pvoff=-6.301879797e-14 nfactor='1.338486025e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.854252010e-05 wnfactor=-3.859840068e-09 pnfactor=7.715384133e-14 eta0=0.08 etab=-0.07 u0=2.128410307e-02 lu0=-2.074325610e-07 wu0=-5.732509211e-09 pu0=1.145863814e-13 ua=1.368212397e-09 lua=-4.335209226e-14 wua=-1.330909162e-15 pua=2.660337022e-20 ub=1.679787904e-19 lub=2.487685152e-23 wub=8.973976729e-25 pub=-1.793796542e-29 uc=-1.117224743e-10 luc=1.211222431e-16 wuc=4.137206980e-18 puc=-8.269809248e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.421845430e+05 lvsat=-1.239880483e+00 wvsat=-2.888185426e-02 pvsat=5.773156301e-7 a0=2.078607149e+00 la0=-1.228530240e-05 wa0=-2.651577759e-07 pa0=5.300204312e-12 ags=1.426154198e-01 lags=-5.861820045e-07 wags=-1.749214772e-08 pags=3.496482668e-13 a1=0.0 a2=1.522317962e+00 la2=-1.104021193e-05 wa2=-2.571713939e-07 pa2=5.140565560e-12 b0=-3.095236262e-07 lb0=4.142166124e-12 wb0=5.125425880e-14 pb0=-1.024514716e-18 b1=-7.552324297e-09 lb1=1.496792631e-13 wb1=3.686839358e-15 pb1=-7.369575264e-20 keta=7.873486781e-02 lketa=-1.106855868e-06 wketa=-2.610002932e-08 pketa=5.217100931e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-3.880260953e-01 lpclm=8.056036225e-06 wpclm=1.869131312e-07 ppclm=-3.736182281e-12 pdiblc1=0.39 pdiblc2=9.024796093e-03 lpdiblc2=-1.548665147e-07 wpdiblc2=-4.168393459e-09 ppdiblc2=8.332147496e-14 pdiblcb=-0.225 drout=0.56 pscbe1=4.384806970e+08 lpscbe1=7.226362351e+03 wpscbe1=2.117136573e+02 ppscbe1=-4.231916773e-3 pscbe2=3.320298000e-09 lpscbe2=1.347315202e-13 wpscbe2=3.247657028e-15 ppscbe2=-6.491699414e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-3.248929186e-10 lalpha0=6.494242313e-15 walpha0=1.512772905e-16 palpha0=-3.023862094e-21 alpha1=-3.248929186e-10 lalpha1=6.494242313e-15 walpha1=1.512772905e-16 palpha1=-3.023862094e-21 beta0=1.177210880e+02 lbeta0=-1.753445424e-03 wbeta0=-4.084486844e-05 pbeta0=8.164427654e-10 agidl=3.536648616e-09 lagidl=-3.350594789e-14 wagidl=-5.676323615e-16 pagidl=1.134632948e-20 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.432067107e-01 lkt1=4.096853045e-06 wkt1=1.164460877e-07 pkt1=-2.327625709e-12 kt2=-7.467703956e-02 lkt2=3.224412527e-07 wkt2=5.553115523e-09 pkt2=-1.110005043e-13 at=-5.657680575e+04 lat=2.549916296e+00 wat=7.830376234e-02 pat=-1.565203726e-6 ute=5.912473887e-01 lute=-1.347704362e-05 wute=-1.854629326e-08 pute=3.707194450e-13 ua1=6.134683819e-09 lua1=-8.084466128e-14 wua1=-1.385827039e-15 pua1=2.770111652e-20 ub1=-5.657513470e-18 lub1=8.852297894e-23 wub1=1.765490015e-24 pub1=-3.529015039e-29 uc1=-1.323423940e-10 luc1=2.049926460e-15 wuc1=2.235391544e-17 puc1=-4.468295096e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.182 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.001192492e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-9.791770030e-08 wvth0=-3.958481478e-08 pvth0=7.784550307e-14 k1=5.348733406e-01 lk1=3.271326537e-08 wk1=-4.364197099e-08 pk1=-5.115496977e-14 k2=2.688621804e-02 lk2=-1.410272908e-07 wk2=-6.736157027e-09 pk2=8.417784970e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.023867703e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=2.156961182e-06 wvoff=1.034093281e-07 pvoff=-8.639560113e-13 nfactor='1.054942708e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.589061313e-05 wnfactor=-7.754151783e-07 pnfactor=6.241009136e-12 eta0=0.08 etab=-0.07 u0=-1.858275187e-02 lu0=1.110585605e-07 wu0=1.604451965e-08 pu0=-5.938747115e-14 ua=-7.304475204e-09 lua=2.593288153e-14 wua=3.780973236e-15 pua=-1.423479372e-20 ub=5.184541336e-18 lub=-1.519981451e-23 wub=-2.418352441e-24 pub=8.551131192e-30 uc=-8.496157175e-11 luc=-9.266712812e-17 wuc=-1.291118286e-17 puc=5.349927763e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-9.958154602e+04 lvsat=6.915573731e-01 wvsat=9.545760975e-02 pvsat=-4.160161837e-7 a0=-2.386114571e-01 la0=6.226655804e-06 wa0=8.247078741e-07 pa0=-3.406590684e-12 ags=-5.369205286e-03 lags=5.960479275e-07 wags=2.971107168e-08 pags=-2.745211655e-14 a1=0.0 a2=-5.174269096e-01 la2=5.255044677e-06 wa2=7.715141817e-07 pa2=-3.077469774e-12 b0=3.155743323e-07 lb0=-8.516602034e-13 wb0=-1.508917569e-13 pb0=5.904035247e-19 b1=-5.011079796e-08 lb1=4.896733765e-13 wb1=2.168927110e-14 pb1=-2.175148395e-19 keta=-9.938390274e-02 lketa=3.161118346e-07 wketa=6.261515623e-08 pketa=-1.870239913e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-7.897111865e-01 lpclm=1.126504620e-05 wpclm=2.246038229e-07 ppclm=-4.037288317e-12 pdiblc1=0.39 pdiblc2=-2.054616505e-02 lpdiblc2=8.137204970e-08 wpdiblc2=1.216857279e-08 ppdiblc2=-4.719242458e-14 pdiblcb=-0.225 drout=0.56 pscbe1=1.884557909e+09 lpscbe1=-4.326160507e+03 wpscbe1=-6.351409718e+02 ppscbe1=2.533494768e-3 pscbe2=3.302779523e-08 lpscbe2=-1.025978132e-13 wpscbe2=-1.078530388e-14 ppscbe2=4.719050623e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=9.746787557e-10 lalpha0=-3.887866848e-15 walpha0=-4.538318716e-16 palpha0=1.810276338e-21 alpha1=9.746787557e-10 lalpha1=-3.887866848e-15 walpha1=-4.538318716e-16 palpha1=1.810276338e-21 beta0=-2.331632640e+02 lbeta0=1.049724049e-03 wbeta0=1.225346053e-04 pbeta0=-4.887746111e-10 agidl=2.248815107e-09 lagidl=-2.321761340e-14 wagidl=-1.063345388e-15 pagidl=1.530651641e-20 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=2.832074918e-01 lkt1=-3.304149585e-06 wkt1=-4.082542109e-07 pkt1=1.864136765e-12 kt2=-1.015288132e-02 lkt2=-1.930338593e-07 wkt2=-1.665934657e-08 pkt2=6.645196775e-14 at=3.076922906e+05 lat=-3.601821589e-01 wat=-1.669313473e-01 pat=3.939476842e-7 ute=-1.773777213e+00 lute=5.416830465e-06 wute=-8.032099971e-08 pute=8.642295441e-13 ua1=-1.004325146e-08 lua1=4.839876052e-14 wua1=4.157481117e-15 pua1=-1.658365170e-20 ub1=1.195721866e-17 lub1=-5.219882614e-23 wub1=-5.296470045e-24 pub1=2.112693047e-29 uc1=2.167821799e-09 luc1=-1.632578625e-14 wuc1=-9.470643324e-16 puc1=7.297726848e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.183 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.058229668e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.295961803e-07 wvth0=-3.077960458e-09 pvth0=-6.777559292e-14 k1=4.420413699e-01 lk1=4.030079283e-07 wk1=-3.259001331e-08 pk1=-9.523979222e-14 k2=1.244243493e-02 lk2=-8.341291769e-08 wk2=1.471276377e-08 pk2=-1.379106991e-15 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.583304515e-01 ldsub=-1.190001388e-06 wdsub=2.259675247e-14 pdsub=-9.013550883e-20 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.782022527e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.185143643e-07 wvoff=-2.051935382e-07 pvoff=3.670207040e-13 nfactor='6.240287060e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.297986226e-06 wnfactor=1.373411130e-06 pnfactor=-2.330379661e-12 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391132325e-01 letab=2.756836997e-7 u0=1.327827155e-02 lu0=-1.603091998e-08 wu0=-1.159826716e-09 pu0=9.238429931e-15 ua=-3.069262731e-09 lua=9.039169554e-15 wua=1.566218255e-15 pua=-5.400424015e-21 ub=6.031517940e-18 lub=-1.857829408e-23 wub=-3.002336697e-24 pub=1.088056847e-29 uc=-8.830803216e-11 luc=-7.931853261e-17 wuc=-2.638083478e-17 puc=1.072279681e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.787700283e+05 lvsat=-4.187508712e-01 wvsat=-5.581668455e-02 pvsat=1.873973106e-7 a0=1.823564999e+00 la0=-1.999097994e-06 wa0=-2.488887635e-07 pa0=8.758467362e-13 ags=-6.119319565e-01 lags=3.015547889e-06 wags=3.346854552e-07 pags=-1.243955286e-12 a1=0.0 a2=0.8 b0=-1.463333337e-07 lb0=9.908294282e-13 wb0=1.317094878e-13 pb0=-5.368561022e-19 b1=1.203930770e-07 lb1=-1.904444152e-13 wb1=-5.447609155e-14 pb1=8.629889059e-20 keta=2.476080193e-04 lketa=-8.130530974e-08 wketa=1.305224933e-08 pketa=1.067600116e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=2.759158628e+00 lpclm=-2.890934136e-06 wpclm=-1.260104079e-06 ppclm=1.885018491e-12 pdiblc1=0.39 pdiblc2=-7.745269496e-04 lpdiblc2=2.505555624e-09 wpdiblc2=6.988029947e-10 ppdiblc2=-1.441003946e-15 pdiblcb=-1.195605023e+00 lpdiblcb=3.871617257e-06 wpdiblcb=4.519350518e-07 ppdiblcb=-1.802710170e-12 drout=0.56 pscbe1=800000000.0 pscbe2=4.818903939e-09 lpscbe2=9.923786967e-15 wpscbe2=2.283964872e-15 ppscbe2=-4.941107795e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-9.944350000e-11 lalpha0=3.966671938e-16 alpha1=-9.944350000e-11 lalpha1=3.966671938e-16 beta0=5.062987286e+01 lbeta0=-8.228988095e-05 wbeta0=2.147046717e-06 pbeta0=-8.564290239e-12 agidl=-5.026033247e-09 lagidl=5.800810955e-15 wagidl=3.471259158e-15 pagidl=-2.781431627e-21 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-9.578050196e-01 lkt1=1.646087992e-06 wkt1=3.057690869e-07 pkt1=-9.840093464e-13 kt2=-5.655244364e-02 lkt2=-7.952037149e-09 wkt2=-3.852746317e-09 pkt2=1.536810420e-14 at=2.778422636e+05 lat=-2.411142819e-01 wat=-6.807471536e-02 pat=-3.785691357e-10 ute=-3.615564910e+00 lute=1.276348216e-05 wute=2.062825386e-06 pute=-7.684502778e-12 ua1=-3.949854351e-10 lua1=9.913081626e-15 wua1=1.913990138e-15 pua1=-7.634657842e-21 ub1=-1.544915052e-18 lub1=1.659429959e-24 wub1=-2.029866285e-25 pub1=8.096872730e-31 uc1=-3.810527422e-09 luc1=7.521071603e-15 wuc1=1.722458408e-15 puc1=-3.350652326e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.184 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.039417136e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=9.218050111e-08 wvth0=-2.436597837e-08 pvth0=-2.543649272e-14 k1=6.750746429e-01 lk1=-6.046495744e-08 wk1=-9.872576197e-08 pk1=3.629561422e-14 k2=-2.822260898e-02 lk2=-2.535431808e-09 wk2=1.345277469e-08 pk2=1.126847487e-15 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=3.099377798e+00 ldsub=-5.647153224e-06 wdsub=-1.662802093e-06 pdsub=3.307097154e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-7.736374448e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.679548262e-07 wvoff=5.163084717e-08 pvoff=-1.437696114e-13 nfactor='9.018681866e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.227879852e-06 wnfactor=-6.114842963e-07 pnfactor=1.617319306e-12 eta0=-1.519541026e+00 leta0=3.023163996e-06 weta0=6.066980445e-07 peta0=-1.206643540e-12 etab=-3.242478655e+00 letab=6.447874088e-06 wetab=1.899006599e-06 petab=-3.776877255e-12 u0=7.323988927e-03 lu0=-4.188625908e-09 wu0=3.192694080e-09 pu0=5.818318953e-16 ua=1.219224695e-09 lua=5.099255679e-16 wua=-8.772250411e-16 pua=-5.407329460e-22 ub=-2.684319370e-18 lub=-1.243626726e-24 wub=2.060338836e-24 pub=8.115649823e-31 uc=-2.517262462e-10 luc=2.456990507e-16 wuc=7.811128004e-17 puc=-1.005932643e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.587901898e+05 lvsat=2.526125199e-01 wvsat=1.023597558e-01 pvsat=-1.271950663e-7 a0=-1.052230102e-01 la0=1.837010613e-06 wa0=6.676304502e-07 pa0=-9.469908324e-13 ags=2.157354643e+00 lags=-2.492203149e-06 wags=-1.115236789e-06 pags=1.639751569e-12 a1=0.0 a2=0.8 b0=4.950739142e-07 lb0=-2.848462048e-13 wb0=-2.159724499e-13 pb0=1.546380732e-19 b1=4.275237513e-07 lb1=-8.012873994e-13 wb1=-2.445647166e-13 pb1=4.643604542e-19 keta=-1.290819922e-01 lketa=1.759144522e-07 wketa=6.550315553e-08 pketa=-9.364203266e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.107973809e+00 lpclm=3.930578153e-07 wpclm=-1.130567811e-07 ppclm=-3.963094679e-13 pdiblc1=4.121363472e-01 lpdiblc1=-4.402631691e-08 wpdiblc1=-9.685305112e-09 ppdiblc1=1.926281278e-14 pdiblc2=5.399081098e-04 lpdiblc2=-1.086848325e-10 wpdiblc2=-5.117563388e-11 ppdiblc2=5.060604908e-17 pdiblcb=1.716210045e+00 lpdiblcb=-1.919604377e-06 wpdiblcb=-9.038701037e-07 ppdiblcb=8.938100294e-13 drout=8.015169287e-01 ldrout=-4.803457740e-07 wdrout=-2.435715807e-07 pdrout=4.844322098e-13 pscbe1=800000000.0 pscbe2=1.015329920e-08 lpscbe2=-6.856317339e-16 wpscbe2=-2.307566904e-16 ppscbe2=6.034647795e-23 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.134202365e-11 lalpha0=1.763291894e-16 walpha0=5.192006143e-17 palpha0=-1.032622526e-22 alpha1=-6.673993786e-10 lalpha1=1.526257602e-15 walpha1=4.494059589e-16 palpha1=-8.938100294e-22 beta0=1.119916002e+01 lbeta0=-3.867319100e-06 wbeta0=-3.820958616e-06 pbeta0=3.305296529e-12 agidl=2.875600971e-09 lagidl=-9.914512293e-15 wagidl=-1.087769216e-15 pagidl=6.285883135e-21 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=2.763963195e-01 lkt1=-8.085780255e-07 wkt1=-4.119049211e-07 pkt1=4.433509579e-13 kt2=-8.325143714e-02 lkt2=4.514879005e-08 wkt2=1.405519212e-08 pkt2=-2.024845732e-14 at=2.142530865e+05 lat=-1.146436752e-01 wat=-1.088087953e-01 pat=8.063622035e-8 ute=6.757041188e+00 lute=-7.866282934e-06 wute=-3.668456273e-06 pute=3.714271374e-12 ua1=8.872030529e-09 lua1=-8.517808414e-15 wua1=-3.429118983e-15 pua1=2.992091596e-21 ub1=-1.093224513e-18 lub1=7.610761966e-25 wub1=-2.764821611e-25 pub1=9.558603327e-31 uc1=3.050590158e-11 luc1=-1.182443435e-16 wuc1=-1.523980640e-17 puc1=1.054035220e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.185 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.574509176e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.112656630e-08 wvth0=-5.680063883e-08 pvth0=6.637169963e-15 k1=1.036233135e+00 lk1=-4.176037558e-07 wk1=-2.674904405e-07 pk1=2.031819418e-13 k2=-2.039832981e-01 lk2=1.712690408e-07 wk2=9.838001200e-08 pk2=-8.285514968e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-8.949702736e+00 ldsub=6.267821044e-06 wdsub=4.969690856e-06 pdsub=-3.251576149e-12 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.532764546e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.772754614e-08 wvoff=-1.435737810e-07 pvoff=4.926238927e-14 nfactor='6.489687589e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.727033282e-06 wnfactor=1.224409451e-06 pnfactor=-1.981409442e-13 eta0=4.861051927e+00 leta0=-3.286412958e-06 weta0=-2.283895339e-06 peta0=1.651777539e-12 etab=6.487716274e+00 letab=-3.174023772e-06 wetab=-3.800221049e-06 petab=1.858917989e-12 u0=-6.421932875e-02 lu0=6.655841464e-08 wu0=3.529326447e-08 pu0=-3.116145915e-14 ua=-6.591124033e-09 lua=8.233345115e-15 wua=2.363224143e-15 pua=-3.745115931e-21 ub=-8.487567513e-18 lub=4.495031265e-24 wub=5.066304269e-24 pub=-2.160944055e-30 uc=1.576238271e-10 luc=-1.590949563e-16 wuc=-1.151140133e-16 puc=9.048143153e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.425073055e+05 lvsat=-4.533153438e-02 wvsat=-5.376875336e-02 pvsat=2.719573252e-8 a0=1.344493545e+00 la0=4.034294024e-07 wa0=3.073766263e-08 pa0=-3.171866615e-13 ags=-1.939894728e+00 lags=1.559443836e-06 wags=1.073854730e-06 pags=-5.249753618e-13 a1=0.0 a2=2.913840811e+00 la2=-2.090313763e-06 wa2=-1.061644519e-06 pa2=1.049828416e-12 b0=4.094350734e-07 lb0=-2.001605243e-13 wb0=-1.178612068e-13 pb0=5.761880816e-20 b1=-7.570439749e-07 lb1=3.700960880e-13 wb1=4.450354859e-13 pb1=-2.175644980e-19 keta=1.935815657e-01 lketa=-1.431578603e-07 wketa=-8.964129099e-08 pketa=5.977565617e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.061344774e+00 lpclm=4.391678689e-07 wpclm=-1.417790393e-07 ppclm=-3.679068884e-13 pdiblc1=4.431003231e-01 lpdiblc1=-7.464566375e-08 wpdiblc1=1.456474821e-07 ppdiblc1=-1.343411205e-13 pdiblc2=-2.882175809e-03 lpdiblc2=3.275311292e-09 wpdiblc2=1.725747505e-09 ppdiblc2=-1.706539935e-15 pdiblcb=2.488695745e-01 lpdiblcb=-4.685954062e-07 wpdiblcb=-2.775084480e-07 ppdiblcb=2.744197790e-13 drout=1.975396214e+00 ldrout=-1.641159782e-06 wdrout=-5.971208369e-07 pdrout=8.340464627e-13 pscbe1=3.957407796e+09 lpscbe1=-3.122265847e+03 wpscbe1=-1.470158533e+03 ppscbe1=1.453795668e-3 pscbe2=-3.195998947e-07 lpscbe2=3.253974091e-13 wpscbe2=1.530238043e-13 ppscbe2=-1.514884912e-19 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=2.773159527e-10 lalpha0=-8.668444980e-17 walpha0=-1.038401229e-16 palpha0=5.076432086e-23 alpha1=1.634798757e-09 lalpha1=-7.503170684e-16 walpha1=-8.988119177e-16 palpha1=4.394021822e-22 beta0=5.113065223e+00 lbeta0=2.151037458e-06 wbeta0=-3.330506028e-07 pbeta0=-1.437910686e-13 agidl=-8.023447427e-09 lagidl=8.632296966e-16 wagidl=5.781596156e-15 pagidl=-5.070262000e-22 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.732833718e-01 lkt1=1.305317309e-07 wkt1=1.164958543e-07 pkt1=-7.916871696e-14 kt2=-1.613356663e-02 lkt2=-2.122205856e-08 wkt2=-1.269939897e-08 pkt2=6.208355176e-15 at=1.162303488e+05 lat=-1.771193063e-02 wat=-5.392306603e-02 pat=2.636136929e-8 ute=-1.870039733e+00 lute=6.647785763e-07 wute=1.776831840e-08 pute=6.907446245e-14 ua1=-2.421503566e-09 lua1=2.650028647e-15 wua1=-3.411093850e-17 pua1=-3.651300094e-22 ub1=4.668020406e-19 lub1=-7.815872610e-25 wub1=1.212877246e-24 pub1=-5.169225039e-31 uc1=-1.103061339e-10 luc1=2.100045407e-17 wuc1=1.806666692e-16 puc1=-8.832251459e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.186 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.214828160e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-6.457159531e-09 wvth0=-3.398312060e-08 pvth0=-4.517630174e-15 k1=8.188028463e-01 lk1=-3.113086104e-07 wk1=-3.047637114e-07 pk1=2.214037258e-13 k2=-1.553872427e-01 lk2=1.475118872e-07 wk2=1.268195278e-07 pk2=-9.675837577e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=6.366663739e+00 ldsub=-1.219891035e-06 wdsub=-3.022304140e-06 pdsub=6.554704447e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-5.902739157e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=6.813340268e-08 wvoff=-1.754827063e-08 pvoff=-1.234770198e-14 nfactor='-8.624535878e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=5.661857144e-06 wnfactor=7.567397592e-06 pnfactor=-3.299037557e-12 eta0=-4.108147213e+00 leta0=1.098359425e-06 weta0=2.140998501e-06 peta0=-5.114203123e-13 etab=-9.184020961e-03 letab=2.115875312e-09 wetab=4.273372071e-09 petab=-9.851980944e-16 u0=1.228863216e-01 lu0=-2.491192465e-08 wu0=-4.967874727e-08 pu0=1.037880823e-14 ua=1.904840340e-08 lua=-4.301050663e-15 wua=-9.180321284e-15 pua=1.898177122e-21 ub=5.498519906e-19 lub=7.690799229e-26 wub=7.966673929e-25 pub=-7.364667538e-32 uc=-3.225775581e-10 luc=7.566109490e-17 wuc=1.341133172e-16 puc=-3.135833352e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.699482999e+04 lvsat=1.361649543e-03 wvsat=-1.025558157e-02 pvsat=5.923448227e-9 a0=5.696410685e+00 la0=-1.724092330e-06 wa0=-2.404335403e-06 pa0=8.732475082e-13 ags=5.810000578e-02 lags=5.826841502e-07 wags=5.549748591e-07 pags=-2.713105594e-13 a1=0.0 a2=-4.697481834e+00 la2=1.630633538e-06 wa2=2.869137901e-06 pa2=-8.718131861e-13 b0=0.0 b1=0.0 keta=-1.510404719e-01 lketa=2.531751523e-08 wketa=5.632197244e-08 pketa=-1.158140442e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=3.925681103e+00 lpclm=-9.611202324e-07 wpclm=-2.160216954e-06 ppclm=6.188468548e-13 pdiblc1=-6.227259153e-01 lpdiblc1=4.464048094e-07 wpdiblc1=2.182871636e-07 ppdiblc1=-1.698524816e-13 pdiblc2=-7.707258018e-03 lpdiblc2=5.634149232e-09 wpdiblc2=6.348467793e-10 ppdiblc2=-1.173231298e-15 pdiblcb=-8.788827743e-01 lpdiblcb=8.272888460e-08 wpdiblcb=4.181909030e-07 ppdiblcb=-6.568676277e-14 drout=-1.466578777e+00 ldrout=4.151853117e-08 wdrout=1.149336726e-06 pdrout=-1.974424604e-14 pscbe1=-5.514807670e+09 lpscbe1=1.508416128e+03 wpscbe1=2.940327369e+03 ppscbe1=-7.023585744e-4 pscbe2=6.699202243e-07 lpscbe2=-1.583492914e-13 wpscbe2=-3.077454202e-13 ppscbe2=7.376775954e-20 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.073916704e+01 lbeta0=-5.993949375e-07 wbeta0=-1.606972851e-06 pbeta0=4.789913008e-13 agidl=-1.223677219e-08 lagidl=2.922997772e-15 wagidl=9.277690851e-15 pagidl=-2.216162014e-21 bgidl=-1.179124819e+08 lbgidl=5.465138750e+02 wbgidl=5.205246456e+02 pbgidl=-2.544688835e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-1.943688208e+00 lkt1=7.515945432e-07 wkt1=6.979518971e-07 pkt1=-3.634251326e-13 kt2=-2.712052184e-02 lkt2=-1.585086577e-08 wkt2=-2.275412971e-08 pkt2=1.112381139e-14 at=2.293166184e+05 lat=-7.299641525e-02 wat=-8.066565581e-02 pat=3.943501915e-8 ute=1.318134179e+00 lute=-8.938240039e-07 wute=-5.781723559e-07 pute=3.604119799e-13 ua1=5.576685961e-09 lua1=-1.260046268e-15 wua1=-1.523518861e-15 pua1=3.629968418e-22 ub1=-1.221665322e-18 lub1=4.385377850e-26 wub1=-1.820449962e-25 pub1=1.650131326e-31 uc1=1.084614330e-10 luc1=-8.594844639e-17 wuc1=-8.587146652e-17 puc1=4.197998384e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.187 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.706050418e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.858193335e-07 wvth0=-4.151075810e-07 pvth0=8.652156968e-14 k1=-6.298412839e+00 lk1=1.388780700e-06 wk1=3.329223700e-06 pk1=-6.466468472e-13 k2=2.782500184e+00 lk2=-5.542612823e-07 wk2=-1.358652162e-06 pk2=2.580762468e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=5.387487042e+00 ldsub=-9.859950972e-07 wdsub=-2.200227547e-06 pdsub=4.591010091e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-1.674265933e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.270665759e-07 wvoff=5.683004807e-07 pvoff=-1.522893932e-13 nfactor='4.507843422e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.166171323e-06 wnfactor=-2.021241812e-05 pnfactor=3.336727024e-12 eta0=4.900000037e-01 leta0=-2.509388253e-16 weta0=-1.704107522e-15 peta0=1.168426467e-22 etab=8.855911077e-03 letab=-2.193323254e-09 wetab=-4.126417165e-09 petab=1.021259560e-15 u0=6.673711861e-02 lu0=-1.149956453e-08 wu0=-2.864488786e-08 pu0=5.354450235e-15 ua=1.238063328e-08 lua=-2.708320415e-15 wua=-6.513081556e-15 pua=1.261053568e-21 ub=-3.346776898e-18 lub=1.007695735e-24 wub=2.452625144e-24 pub=-4.692053034e-31 uc=1.394789572e-10 luc=-3.471034490e-17 wuc=-6.482432146e-17 puc=1.616190021e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.352410285e+05 lvsat=-6.749171990e-02 wvsat=-1.170173406e-01 pvsat=3.142562960e-8 a0=-4.600347823e+00 la0=7.354943751e-07 wa0=2.685085077e-06 pa0=-3.424623619e-13 ags=5.506785593e+00 lags=-7.188433760e-07 wags=-1.982053021e-06 pags=3.347092904e-13 a1=0.0 a2=2.686163724e+00 la2=-1.330978760e-07 wa2=-1.040044856e-06 pa2=6.197329922e-14 b0=0.0 b1=0.0 keta=-2.700592797e-01 lketa=5.374753786e-08 wketa=1.126062763e-07 pketa=-2.502603607e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=9.549166851e-02 lpclm=-4.620288215e-08 wpclm=3.404477442e-07 ppclm=2.151307839e-14 pdiblc1=1.829534444e+00 lpdiblc1=-1.393666226e-07 wpdiblc1=-7.644425520e-07 ppdiblc1=6.489216557e-14 pdiblc2=1.022867181e-01 lpdiblc2=-2.064011184e-08 wpdiblc2=-4.450988237e-08 ppdiblc2=9.610490155e-15 pdiblcb=9.486856462e+00 lpdiblcb=-2.393335247e-06 wpdiblcb=-4.522054030e-06 ppdiblcb=1.114389544e-12 drout=-6.841647336e+00 ldrout=1.325461158e-06 wdrout=3.650360836e-06 pdrout=-6.171638752e-13 pscbe1=7.996773148e+08 lpscbe1=7.509940378e-02 wpscbe1=1.356055240e-01 ppscbe1=-3.496793459e-8 pscbe2=5.045485777e-08 lpscbe2=-1.037759935e-14 wpscbe2=-1.915446704e-14 ppscbe2=4.832038563e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=1.477571885e+01 lbeta0=-1.563606069e-06 wbeta0=-2.649624018e-06 pbeta0=7.280493850e-13 agidl=-1.218911605e-08 lagidl=2.911614151e-15 wagidl=5.675520595e-15 pagidl=-1.355711604e-21 bgidl=4.992544064e+09 lbgidl=-6.742208802e+02 wbgidl=-1.859016352e+03 pbgidl=3.139320747e-4 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=7.845529920e+00 lkt1=-1.586755991e-06 wkt1=-3.916497932e-06 pkt1=7.388284981e-13 kt2=-1.173440897e-01 lkt2=5.700837883e-09 wkt2=3.492681360e-08 pkt2=-2.654435537e-15 at=5.077620567e+05 lat=-1.395086771e-01 wat=-1.875157839e-01 pat=6.495830924e-8 ute=-6.560091088e+00 lute=9.880476656e-07 wute=2.856619414e-06 pute=-4.600567301e-13 ua1=-3.452041285e-10 lua1=1.545156182e-16 wua1=2.973155380e-16 pua1=-7.194587116e-23 ub1=-1.690910674e-18 lub1=1.559424157e-25 wub1=8.127360648e-25 pub1=-7.261021949e-32 uc1=-1.058809044e-09 luc1=1.928774524e-16 wuc1=4.658427252e-16 puc1=-8.980798513e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.188 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='-1.977238765e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.312734016e-07 wvth0=4.289966288e-07 pvth0=-6.166202659e-14 k1=5.014142124e+00 lk1=-5.740765128e-07 wk1=-2.229347261e-06 pk1=3.214273464e-13 k2=-1.617295902e+00 lk2=2.077318020e-07 wk2=8.393207775e-07 pk2=-1.244806661e-13 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-5.070246770e-01 ldsub=1.035850396e-08 wdsub=9.683496291e-07 pdsub=-8.362512053e-14 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='4.858351638e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=-8.542255367e-07 wvoff=-2.775498456e-06 pvoff=4.538916709e-13 nfactor='5.391786822e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-9.530569323e-06 wnfactor=-2.594275507e-05 pnfactor=4.737730238e-12 eta0=7.745943584e+00 leta0=-1.348662234e-06 weta0=-3.378526964e-06 peta0=6.279668065e-13 etab=3.959197557e-01 letab=-7.435768005e-08 wetab=-1.828549683e-07 petab=3.434434469e-14 u0=1.348367508e-02 lu0=-2.758998410e-09 wu0=-4.793375176e-09 pu0=1.460197547e-15 ua=-1.164721104e-09 lua=-4.632897192e-16 wua=-3.095434695e-16 pua=2.349511397e-22 ub=2.280736421e-18 lub=6.315371116e-26 wub=-4.418928819e-25 pub=2.156426123e-32 uc=-7.672994775e-10 luc=1.303383017e-16 wuc=4.043708594e-16 puc=-6.942040324e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.755283976e+05 lvsat=1.135856590e-01 wvsat=4.176558073e-01 pvsat=-6.479047685e-8 a0=-6.935358078e+00 la0=1.243544328e-06 wa0=4.162627355e-06 pa0=-6.515685413e-13 ags=1.250000270e+00 lags=-4.235737183e-14 wags=-1.255811632e-13 pags=1.972252406e-20 a1=0.0 a2=7.693463499e-01 la2=2.097821188e-07 wa2=-5.869303230e-07 pa2=-1.600829949e-14 b0=0.0 b1=0.0 keta=-9.988449067e-01 lketa=1.946176415e-07 wketa=4.253777128e-07 pketa=-8.568021286e-14 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-4.285013399e+00 lpclm=7.633503896e-07 wpclm=2.869001892e-06 ppclm=-4.463035776e-13 pdiblc1=5.165122340e+00 lpdiblc1=-7.733822648e-07 wpdiblc1=-2.258240345e-06 ppdiblc1=3.490770007e-13 pdiblc2=-1.049004960e-01 lpdiblc2=1.579195305e-08 wpdiblc2=5.919108705e-08 ppdiblc2=-8.696929121e-15 pdiblcb=-3.668849702e+01 lpdiblcb=5.948342671e-06 wpdiblcb=1.765861111e-05 ppdiblcb=-2.896146032e-12 drout=1.045574033e+00 ldrout=-7.103624891e-09 wdrout=-2.668906125e-08 pdrout=4.160024129e-15 pscbe1=1.259780903e+09 lpscbe1=-8.543679443e+01 wpscbe1=-2.141737918e+02 ppscbe1=3.979519955e-5 pscbe2=-1.104974066e-07 lpscbe2=1.849389388e-14 wpscbe2=5.541536989e-14 ppscbe2=-8.541819795e-21 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=-7.893512919e-02 lbeta0=1.040021567e-06 wbeta0=5.968381082e-06 pbeta0=-8.004871074e-13 agidl=3.130442945e-08 lagidl=-4.879421419e-15 wagidl=-1.457603105e-14 pagidl=2.271965960e-21 bgidl=1.000001312e+09 lbgidl=-2.042606182e-04 wbgidl=-6.108383255e-04 pbgidl=9.510823774e-11 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.447415107e+00 lkt1=3.525263183e-07 wkt1=1.686375233e-06 pkt1=-2.282002975e-13 kt2=7.944095580e-01 lkt2=-1.631929141e-07 wkt2=-3.740163109e-07 pkt2=7.308860324e-14 at=-2.609334921e+06 lat=4.258219176e-01 wat=1.428116186e+00 pat=-2.287999070e-7 ute=-3.545751960e+00 lute=5.272383744e-07 wute=8.196532909e-07 pute=-1.277593586e-13 ua1=1.536643681e-09 lua1=-1.797084777e-16 wua1=-1.910596230e-15 pua1=3.311959592e-22 ub1=-1.057100144e-18 lub1=5.383464358e-26 wub1=2.172518994e-24 pub1=-3.326626819e-31 uc1=-4.085983784e-11 luc1=2.308804341e-17 wuc1=5.102270534e-17 puc1=-2.174628191e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.189 pmos lmin=2.0e-05 lmax=0.0001 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.0909497+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.43165561 k2=0.019248026 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=3.2465718e-7 voff='-1.02249072+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='11.4566612+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.08 etab=-0.07 u0=0.0109067 ua=-8.0059916e-10 ub=1.41251395e-18 uc=-1.0566299e-10 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.464 ags=0.11329 a1=0.0 a2=0.97 b0=-1.023e-7 b1=-6.41939999999979e-11 keta=0.023361259 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.015 pdiblc1=0.39 pdiblc2=0.0012771588 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=1.0060625e-8 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=1.8604184e-9 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.43825 kt2=-0.058546 at=70990.0 ute=-0.08298 ua1=2.0902e-9 ub1=-1.2289e-18 uc1=-2.9789e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.190 pmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.099879193e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.784904721e-7 k1=4.317673477e-01 lk1=-2.233509594e-9 k2=2.048102620e-02 lk2=-2.464628068e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=-6.116597486e-06 lcit=1.287534022e-10 wcit=-1.482307658e-27 pcit=-2.032879073e-32 voff='-1.194549843e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.439267434e-6 nfactor='1.337657060e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.837681950e-5 eta0=0.08 etab=-0.07 u0=8.972594573e-03 lu0=3.866058195e-8 ua=-1.490134421e-09 lua=1.378303069e-14 ub=2.095288224e-18 lub=-1.364788619e-23 uc=-1.028371403e-10 luc=-5.648554281e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80156.0 a0=1.509137115e+00 la0=-9.022399339e-07 wa0=-8.881784197e-22 ags=1.050481491e-01 lags=1.647452859e-7 a1=0.0 a2=0.97 b0=-1.994466564e-07 lb0=1.941851886e-12 b1=3.657709778e-10 lb1=-8.594514046e-15 wb1=-5.169878828e-32 pb1=-1.240770919e-36 keta=2.268075241e-02 lketa=1.360255782e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.340066551e-02 lpclm=3.196888926e-8 pdiblc1=0.39 pdiblc2=7.248400546e-05 lpdiblc2=2.408008786e-8 pdiblcb=-0.225 drout=0.56 pscbe1=8.931706757e+08 lpscbe1=-1.862376525e+3 pscbe2=1.029517683e-08 lpscbe2=-4.688425941e-15 wpscbe2=6.617444900e-30 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=2.317564549e-09 lagidl=-9.137834950e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.931195419e-01 lkt1=-9.021068602e-7 kt2=-6.275080858e-02 lkt2=8.404937201e-8 at=1.115934318e+05 lat=-8.116167193e-1 ute=5.514161667e-01 lute=-1.268086250e-05 wute=-5.551115123e-23 ua1=3.158391808e-09 lua1=-2.135194718e-14 pua1=1.323488980e-35 ub1=-1.865832633e-18 lub1=1.273156360e-23 pub1=-6.162975822e-45 uc1=-8.433367566e-11 luc1=1.090286431e-15 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.191 pmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.086207407e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=6.926834990e-8 k1=4.411450137e-01 lk1=-7.715046481e-8 k2=1.241921041e-02 lk2=3.975851759e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.56 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.017791248e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.014732292e-7 nfactor='8.884095162e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.487017214e-6 eta0=0.08 etab=-0.07 u0=1.587549891e-02 lu0=-1.648582346e-8 ua=8.157880917e-10 lua=-4.638684493e-15 ub=-9.269181748e-21 lub=3.165149325e-24 uc=-1.126904653e-10 luc=2.223138962e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.054294065e+05 lvsat=-2.019059592e-1 a0=1.532584651e+00 la0=-1.089559245e-6 ags=5.844021883e-02 lags=5.370899819e-7 a1=0.0 a2=1.139526975e+00 la2=-1.354328965e-6 b0=-8.490589332e-09 lb0=4.163286904e-13 b1=-3.529512926e-09 lb1=2.252440268e-14 pb1=-3.308722450e-36 keta=3.509246699e-02 lketa=-8.555301647e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-3.073374523e-01 lpclm=2.594304016e-6 pdiblc1=0.39 pdiblc2=5.587850927e-03 lpdiblc2=-1.998146148e-8 pdiblcb=-0.225 drout=0.56 pscbe1=5.204879729e+08 lpscbe1=1.114937140e+3 pscbe2=9.864577265e-09 lpscbe2=-1.248422033e-15 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=0.0 alpha1=0.0 beta0=30.0 agidl=-3.489440034e-11 lagidl=9.655653779e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-5.935857243e-01 lkt1=6.993914107e-7 kt2=-4.593157427e-02 lkt2=-5.031730436e-8 at=-5.082029532e+04 lat=4.858854327e-01 wat=7.275957614e-18 pat=1.164153218e-22 ute=-1.946279800e+00 lute=7.272905874e-6 ua1=-1.114375423e-09 lua1=1.278263477e-14 pua1=1.654361225e-36 ub1=5.821761488e-19 lub1=-6.825260318e-24 pub1=-1.540743956e-45 uc1=1.338450270e-10 luc1=-6.527148612e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.192 pmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.064840095e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.596307788e-8 k1=3.720489440e-01 lk1=1.984647748e-7 k2=4.404052043e-02 lk2=-8.637477729e-8 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=8.583305000e-01 ldsub=-1.190001582e-6 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-8.188892009e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=3.697230987e-7 nfactor='9.189913861e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-3.706888247e-6 eta0=1.590575825e-01 leta0=-3.153504191e-7 etab=-1.391132325e-01 letab=2.756836997e-7 u0=1.078735248e-02 lu0=3.810131197e-9 ua=2.944491542e-10 lua=-2.559131245e-15 ub=-4.164950337e-19 lub=4.789520309e-24 uc=-1.449652236e-10 luc=1.509712047e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.889449718e+04 lvsat=-1.628425534e-2 a0=1.289035351e+00 la0=-1.180727503e-7 ags=1.068602294e-01 lags=3.439488544e-7 a1=0.0 a2=0.8 b0=1.365345028e-07 lb0=-1.621575488e-13 b1=3.396690349e-09 lb1=-5.103321782e-15 keta=2.827946504e-02 lketa=-5.837683738e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=5.287739745e-02 lpclm=1.157453809e-6 pdiblc1=0.39 pdiblc2=7.262676750e-04 lpdiblc2=-5.892378908e-10 pdiblcb=-0.225 drout=0.56 pscbe1=800000000.0 pscbe2=9.724094998e-09 lpscbe2=-6.880565344e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=-9.944350000e-11 lalpha0=3.966671938e-16 alpha1=-9.944350000e-11 lalpha1=3.966671938e-16 beta0=5.524100961e+01 lbeta0=-1.006831060e-4 agidl=2.429068011e-09 lagidl=-1.727719663e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-3.011155013e-01 lkt1=-4.672342876e-7 kt2=-6.482685146e-02 lkt2=2.505349996e-8 at=1.316405906e+05 lat=-2.419273215e-1 ute=8.146926502e-01 lute=-3.740254304e-06 wute=2.220446049e-22 pute=-6.661338148e-28 ua1=3.715623896e-09 lua1=-6.483604617e-15 ub1=-1.980862298e-18 lub1=3.398366850e-24 uc1=-1.112640540e-10 luc1=3.249933986e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.193 pmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-09*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.091747092e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.755143993e-8 k1=4.630447947e-01 lk1=1.748585722e-8 k2=6.694422700e-04 lk2=-1.153410749e-10 wk2=4.336808690e-25 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-4.717638000e-01 ldsub=1.455383069e-06 pdsub=-2.220446049e-28 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.627516895e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.918588626e-8 nfactor='7.705418540e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-7.544200379e-7 eta0=-2.165569650e-01 leta0=4.316980860e-07 weta0=3.035766083e-24 peta0=3.209238431e-29 etab=8.359510565e-01 letab=-1.663592413e-06 wetab=2.190088388e-22 petab=1.899522206e-28 u0=1.418082576e-02 lu0=-2.939046001e-9 ua=-6.647606861e-10 lua=-6.513875702e-16 ub=1.740597915e-18 lub=4.993428553e-25 uc=-8.396939611e-11 luc=2.965843340e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.104425915e+04 lvsat=-2.055985244e-2 a0=1.328623436e+00 la0=-1.968083056e-7 ags=-2.378002026e-01 lags=1.029433648e-06 pags=2.220446049e-28 a1=0.0 a2=0.8 b0=3.123747616e-08 lb0=4.726454853e-14 b1=-9.771929255e-08 lb1=1.960032231e-13 wb1=2.481541838e-29 pb1=3.887748879e-35 keta=1.159683213e-02 lketa=-2.519724925e-08 wketa=2.602085214e-24 pketa=-8.673617380e-31 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=8.651657345e-01 lpclm=-4.580820963e-07 wpclm=-4.440892099e-22 pdiblc1=3.913355579e-01 lpdiblc1=-2.656251107e-9 pdiblc2=0.00043 pdiblcb=-0.225 drout=2.784068077e-01 ldrout=5.600522523e-7 pscbe1=800000000.0 pscbe2=9.657711168e-09 lpscbe2=-5.560277248e-16 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.228489143e-10 lalpha0=-4.544352013e-17 alpha1=2.977740000e-10 lalpha1=-3.933467754e-16 beta0=2.993021526e+00 lbeta0=3.231350053e-6 agidl=5.394372676e-10 lagidl=3.585457931e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-6.082373987e-01 lkt1=1.435912404e-7 kt2=-5.306559515e-02 lkt2=1.661890126e-9 at=-1.943173781e+04 lat=5.853590038e-02 pat=-7.275957614e-24 ute=-1.121573381e+00 lute=1.107271173e-7 ua1=1.507432243e-09 lua1=-2.091798484e-15 pua1=-4.135903063e-37 ub1=-1.687015530e-18 lub1=2.813943829e-24 wub1=1.925929944e-40 pub1=-5.777789833e-46 uc1=-2.224094860e-12 luc1=1.081270951e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.194 pmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.079439653e+00+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.538098290e-8 k1=4.617533202e-01 lk1=1.876295759e-8 k2=7.303995037e-03 lk2=-6.676051270e-09 wk2=4.336808690e-25 pk2=6.505213035e-31 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=1.723527600e+00 ldsub=-7.154747378e-7 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.616248165e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.807155544e-08 wvoff=4.440892099e-22 nfactor='9.119308722e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.152573622e-6 eta0=-4.398980000e-02 leta0=2.610515935e-7 etab=-1.673884872e+00 letab=8.183090420e-7 u0=1.157877459e-02 lu0=-3.659556598e-10 ua=-1.515710622e-09 lua=1.900912925e-16 ub=2.393156055e-18 lub=-1.459523120e-25 uc=-8.960249234e-11 luc=3.522883326e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.703004424e+04 lvsat=1.307578426e-2 a0=1.410507743e+00 la0=-2.777812396e-7 ags=3.663853228e-01 lags=4.319727072e-7 a1=0.0 a2=6.337842000e-01 la2=1.643658181e-7 b0=1.563087032e-07 lb0=-7.641463571e-14 b1=1.987430926e-07 lb1=-9.715953568e-14 keta=1.062116491e-03 lketa=-1.477978500e-8 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=7.568509154e-01 lpclm=-3.509728211e-7 pdiblc1=7.559023000e-01 lpdiblc1=-3.631653654e-7 pdiblc2=8.241514375e-04 lpdiblc2=-3.897645320e-10 pdiblcb=-3.471255631e-01 lpdiblcb=1.207663056e-7 drout=6.929807845e-01 ldrout=1.500924839e-7 pscbe1=800000000.0 pscbe2=9.043950024e-09 lpscbe2=5.090225685e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=5.430217145e-11 lalpha0=2.234029744e-17 alpha1=-2.955480000e-10 lalpha1=1.933715508e-16 beta0=4.397784152e+00 lbeta0=1.842222435e-6 agidl=4.393483380e-09 lagidl=-2.256926483e-16 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.230893210e-01 lkt1=-3.949613924e-8 kt2=-4.340761934e-02 lkt2=-7.888592413e-9 at=4.216756200e+02 lat=3.890345544e-2 ute=-1.831879340e+00 lute=8.131273709e-7 ua1=-2.494762429e-09 lua1=1.865851762e-15 wua1=8.271806126e-31 pua1=-4.135903063e-37 ub1=3.071655861e-18 lub1=-1.891763550e-24 pub1=7.703719778e-46 uc1=2.777053201e-10 luc1=-1.686867054e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.195 pmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-9.944671694e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.615951504e-8 k1=1.642725377e-01 lk1=1.641923878e-7 k2=1.169785987e-01 lk2=-6.029267476e-08 wk2=2.775557562e-23 pk2=6.938893904e-30 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=-1.242326091e-01 ldsub=1.878397956e-07 pdsub=5.551115123e-29 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-6.279617196e-01+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=4.161467724e-8 nfactor='7.627697891e+00+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.423369835e-6 eta0=0.49 etab=-6.25e-6 u0=1.619302260e-02 lu0=-2.621723083e-9 ua=-6.678498755e-10 lua=-2.244023905e-16 ub=2.260826543e-18 lub=-8.126038331e-26 wub=-1.540743956e-39 uc=-3.454710167e-11 luc=8.313904430e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.496927800e+04 lvsat=1.408323105e-2 a0=5.327040663e-01 la0=1.513506437e-7 ags=1.25 a1=0.0 a2=1.464464770e+00 la2=-2.417289920e-7 b0=0.0 b1=0.0 keta=-3.007975172e-02 lketa=4.445401076e-10 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=-7.137409036e-01 lpclm=3.679554014e-07 wpclm=2.775557562e-23 ppclm=5.551115123e-29 pdiblc1=-1.539182482e-01 lpdiblc1=8.161860606e-08 wpdiblc1=-2.775557562e-23 ppdiblc1=-1.040834086e-29 pdiblc2=-6.343819909e-03 lpdiblc2=3.114441620e-09 wpdiblc2=7.318364664e-25 ppdiblc2=-5.624298770e-31 pdiblcb=1.925112622e-02 lpdiblcb=-5.834426652e-8 drout=1.001811303e+00 ldrout=-8.854919108e-10 pscbe1=8.000300498e+08 lpscbe1=-1.469046821e-2 pscbe2=8.986204433e-09 lpscbe2=7.913234404e-17 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=7.287927943e+00 lbeta0=4.293178398e-7 agidl=7.688598287e-09 lagidl=-1.836575473e-15 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-4.447214558e-01 lkt1=-2.892083750e-8 kt2=-7.598876628e-02 lkt2=8.039352891e-9 at=5.607382532e+04 lat=1.169678902e-2 ute=7.641373640e-02 lute=-1.197798653e-07 pute=-2.775557562e-29 ua1=2.304678064e-09 lua1=-4.804507120e-16 ub1=-1.612636960e-18 lub1=3.982466821e-25 uc1=-7.596169672e-11 luc1=4.210489046e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.196 pmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=5.565e-9 vth0='-1.062117+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' k1=0.85164386 k2=-0.1354293 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=0.66213569 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-0.45374697+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' nfactor='1.6689344+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' eta0=0.49 etab=-6.25e-6 u0=0.0052175 ua=-1.607283e-9 ub=1.9206399e-18 uc=2.58041e-13 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=83927.0 a0=1.166315 ags=1.25 a1=0.0 a2=0.45249595 b0=0.0 b1=0.0 keta=-0.028218739 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=0.82665932 pdiblc1=0.18776805 pdiblc2=0.0066944085 pdiblcb=-0.225 drout=0.9981043 pscbe1=799968550.0 pscbe2=9.3174823e-9 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=9.0852145 agidl=0.0 bgidl=1000000000.0 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.4765e-8 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=-0.565795 kt2=-0.042333 at=105041.0 ute=-0.42503 ua1=2.9333e-10 ub1=5.4574e-20 uc1=-5.8335e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.model sky130_fd_pr__pfet_01v8_hvt__model.197 pmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.6e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre*(4.23e-9*0.948*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))' toxm=4.23e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-2.2811e-8 lint=-2.935e-9 vth0='5.074060142e-01+sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.917272426e-07 wvth0=-7.279086425e-07 pvth0=1.352963794e-13 k1=-1.747554175e+00 lk1=4.831129388e-07 wk1=9.190472936e-07 pk1=-1.708233205e-13 k2=-2.219594058e-01 lk2=1.608335076e-08 wk2=1.896214072e-07 pk2=-3.524493096e-14 k3=-13.778 k3b=2.0 w0=0.0 dvt0=4.05 dvt1=0.3 dvt2=0.03 dvt0w=-4.254 dvt1w=1147200.0 dvt2w=-0.00896 dsub=6.670698446e+00 ldsub=-1.116811559e-06 wdsub=-2.373756167e-06 pdsub=4.412100587e-13 minv=0.0 voffl=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 cit=1.0e-5 voff='-3.576606805e+00+sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))' lvoff=5.804459575e-07 wvoff=1.152003764e-06 pvoff=-2.141229396e-13 nfactor='-1.631964868e+01+sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=3.343537937e-06 wnfactor=6.761378024e-06 pnfactor=-1.256737333e-12 eta0=7.745943542e+00 leta0=-1.348662226e-06 weta0=-3.378526944e-06 peta0=6.279668031e-13 etab=4.457253357e-01 letab=-8.284812984e-08 wetab=-2.060455421e-07 petab=3.829768491e-14 u0=3.911196982e-02 lu0=-6.299965106e-09 wu0=-1.672647303e-08 pu0=3.108949542e-15 ua=1.153628828e-08 lua=-2.442995595e-15 wua=-6.223412863e-15 pua=1.156745749e-21 ub=-2.055422691e-18 lub=7.390307538e-25 wub=1.577118196e-24 pub=-2.931389591e-31 uc=-3.828960618e-10 luc=7.121685309e-17 wuc=2.253841722e-16 puc=-4.189215609e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.714324205e+06 lvsat=-3.030419284e-01 wvsat=-6.951121410e-01 pvsat=1.292004937e-7 a0=1.808836105e+00 la0=-1.194253977e-07 wa0=9.113817138e-08 pa0=-1.693985192e-14 ags=1.249999985e+00 lags=2.731505688e-15 wags=6.842682865e-15 pags=-1.271849293e-21 a1=0.0 a2=-8.632484378e+00 la2=1.688625294e-06 wa2=3.790768904e-06 pa2=-7.045902162e-13 b0=0.0 b1=0.0 keta=-1.472423496e+00 lketa=2.684343382e-07 wketa=6.458863228e-07 pketa=-1.200508908e-13 dwg=-5.722e-9 dwb=-1.7864e-8 pclm=1.940062338e+00 lpclm=-2.069482190e-07 wpclm=-2.953032308e-08 ppclm=5.488801151e-15 pdiblc1=9.440897930e-02 lpdiblc1=1.735265047e-08 wpdiblc1=1.027953514e-07 ppdiblc1=-1.910657197e-14 pdiblc2=6.230151542e-02 lpdiblc2=-1.033569296e-08 wpdiblc2=-1.866184791e-08 ppdiblc2=3.468677671e-15 pdiblcb=-9.647124730e+00 lpdiblcb=1.751290324e-06 wpdiblcb=5.067553259e-06 ppdiblcb=-9.419061243e-13 drout=9.882548598e-01 ldrout=1.830715458e-09 wdrout=6.956739185e-15 pdrout=-1.293049223e-21 pscbe1=1.285433399e+09 lpscbe1=-9.023335140e+01 wpscbe1=-2.261181578e+02 ppscbe1=4.202858199e-5 pscbe2=1.576995002e-08 lpscbe2=-1.199320176e-15 wpscbe2=-3.377489220e-15 ppscbe2=6.277739214e-22 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=531.92 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=-0.32348 prwg=0.02 wr=1.0 alpha0=1.0e-10 alpha1=1.0e-10 beta0=2.257026038e+01 lbeta0=-2.506465477e-06 wbeta0=-4.577582627e-06 pbeta0=8.508352829e-13 agidl=0.0 bgidl=1.000000010e+09 lbgidl=-1.901000977e-06 wbgidl=-4.762187958e-06 pbgidl=8.851480484e-13 cgidl=300.0 egidl=0.1 toxref=4.23e-9 dlcig=0.0 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=1.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=6.265e-9 dwc=-3.2175e-8 xpart=0.0 cgso=5.46384e-11 cgdo=5.46384e-11 cgbo=0.0 cgdl=6.920864e-12 cgsl=6.920864e-12 clc=1.0e-7 cle=0.6 cf=1.2e-11 ckappas=0.6 vfbcv=-0.1446893 acde=0.552 moin=14.504 noff=4.0 voffcv=-0.1375 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.88 noia=1.2e+41 noib=2.0e+25 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-6.0e-8 af=1.0 kf=0.0 tnoia=1.5 tnoib=3.5 rnoia=0.577 rnoib=0.37 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=2.17e-5 jsws=8.2e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=12.8 xjbvs=1.0 pbs=0.6587 cjs=0.000672644022 mjs=0.34629 pbsws=0.7418 cjsws=8.60458928e-11 mjsws=0.26859 pbswgs=1.3925 cjswgs=2.299366688e-10 mjswgs=0.70393 tnom=30.0 kt1=3.606711407e+00 lkt1=-7.755437659e-07 wkt1=-1.598181263e-06 pkt1=2.970539513e-13 kt2=1.111362601e+00 lkt2=-2.144374014e-07 wkt2=-5.215966208e-07 pkt2=9.694916391e-14 at=-1.175221209e+04 lat=2.170835433e-02 wat=2.186245303e-01 pat=-4.063574145e-8 ute=-1.785411394e+00 lute=2.528540896e-07 wute=-4.483453608e-15 pute=8.333396195e-22 ua1=-3.768870207e-11 lua1=6.152644615e-17 wua1=-1.177552437e-15 pua1=2.188716715e-22 ub1=4.060735096e-18 lub1=-7.446251629e-25 wub1=-2.104576860e-25 pub1=3.911777010e-32 uc1=-9.759609062e-10 luc1=1.705591272e-16 wuc1=4.864263350e-16 puc1=-9.041206288e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2556 tpb=0.0019551 tcj=0.0012407 tpbsw=0.00014242 tcjsw=0.0 tpbswg=0.0 tcjswg=2.0e-12 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=2.65e-8 lkvth0=0.0 wkvth0=2.5e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=4.5e-8 lku0=0.0 wku0=2.5e-7 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.4 steta0=0.0
.ends sky130_fd_pr__pfet_01v8_hvt