* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_cm04w5p00l0p25 drain gate source substrate
x0 substrate substrate source substrate sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=150000u
x1 source substrate substrate substrate sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=150000u
x2 drain gate source substrate sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=250000u
x3 source gate drain substrate sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=250000u
x4 drain gate source substrate sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=250000u
x5 source gate drain substrate sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=250000u
.ends