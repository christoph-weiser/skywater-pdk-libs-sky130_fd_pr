* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_g5v0d10v5__toxe_mult=1.042
.param sky130_fd_pr__pfet_g5v0d10v5__rshp_mult=1.0
.param sky130_fd_pr__pfet_g5v0d10v5__overlap_mult=1.1981e+0
.param sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult=1.0559e+0
.param sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult=1.0542e+0
.param sky130_fd_pr__pfet_g5v0d10v5__lint_diff=-1.21275e-8
.param sky130_fd_pr__pfet_g5v0d10v5__wint_diff=2.252e-8
.param sky130_fd_pr__pfet_g5v0d10v5__dlc_diff=-1.21275e-8
.param sky130_fd_pr__pfet_g5v0d10v5__dwc_diff=2.252e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0=-9.7632e-20
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0=6.0196e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0=0.012891
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0=0.38252
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0=-0.0017077
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0=-0.069006
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0=-4769.9
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1=-7.9015e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1=4.1439e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1=-0.02713
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1=0.015985
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1=0.32012
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1=-0.002803
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1=-0.053981
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1=-0.073156
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2=-2.4902e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2=5.9639e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2=0.011096
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2=0.59119
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2=-0.002166
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2=-0.076026
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2=-6616.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3=0.04597
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3=-3.4756e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3=1.367e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3=-6.449e-5
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3=0.0076581
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3=0.34106
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3=-0.0013318
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3=-0.049718
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4=0.44847
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4=-0.0010083
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4=-0.056905
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4=0.016874
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4=-4.2561e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4=3.0864e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4=0.01461
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4=0.0060092
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5=0.0081495
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5=0.51875
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5=-0.0019456
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5=-0.045101
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5=0.016937
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5=-6.3323e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5=9.121e-12
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5=0.010857
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6=0.0073926
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6=0.095219
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6=-0.0016464
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6=-0.051876
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6=-1863.9
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6=-8.2882e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6=2.886e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7=0.014954
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7=0.0095634
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7=-0.053071
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7=0.24848
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7=-0.0012312
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7=-0.01603
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7=-2.7184e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7=4.6643e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8=-0.024268
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8=0.0077753
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8=-0.04579
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8=0.3146
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8=-0.0016667
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8=-0.066818
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8=-3.861e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8=1.2881e-11
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9=0.015574
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9=0.0044227
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9=-0.055474
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9=0.64327
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9=-0.0011345
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9=0.016879
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9=-1.7933e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9=1.5302e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10=0.62279
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10=-0.00099328
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10=-0.045112
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10=0.014396
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10=0.0059166
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10=6.109e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10=-8.7392e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10=0.0055447
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11=13338.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11=0.08928
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11=-0.00022049
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11=-0.11155
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11=0.0053403
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11=8.5687e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11=8.8343e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12=1022.6
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12=0.11878
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12=-0.0019019
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12=-0.05422
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12=0.0034067
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12=4.3051e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12=-4.928e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13=-4.1132e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13=-673.64
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13=-0.044538
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13=-0.0011289
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13=-0.090735
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13=0.0098142
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13=7.0038e-11
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14=4.9102e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14=-2.8249e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14=-0.031865
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14=0.24677
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14=-0.0015275
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14=-0.059832
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14=-0.095284
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14=0.015894
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15=0.012739
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15=6.2456e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15=-1.8609e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15=-6563.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15=0.23246
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15=-0.0017419
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15=-0.070692
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16=-0.050038
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16=-0.048464
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16=0.013921
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16=3.3816e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16=-8.1137e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16=-0.008898
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16=0.30971
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16=-0.0023631
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17=0.011174
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17=-0.0008474
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17=-0.060383
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17=0.00054553
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17=0.0072257
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17=5.2675e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17=-2.9752e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17=0.029451
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18=0.92406
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18=-0.0026389
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18=-0.037376
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18=-0.015684
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18=0.0085502
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18=-1.3071e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18=-9.6709e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18=0.0091247
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19=0.65267
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19=-0.0020078
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19=-0.043644
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19=-0.0047006
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19=0.0073137
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19=3.6802e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19=-6.7659e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19=0.012858
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20=0.06487
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20=-0.00053524
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20=-0.092462
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20=0.011449
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20=6.7256e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20=-1.2735e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20=5702.6
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21=-4825.1
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21=0.13037
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21=-0.0024014
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21=-0.062924
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21=0.014179
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21=4.1947e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21=-9.9157e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22=-0.025754
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22=-0.041992
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22=-0.08788
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22=0.00057436
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22=-0.092463
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22=-0.070061
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22=0.010742
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22=9.382e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22=2.5117e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23=0.0027807
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23=-0.0015768
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23=-0.064703
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23=-0.0054163
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23=0.0087627
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23=1.836e-14
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23=-4.4666e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24=-9.2154e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24=0.01206
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24=0.90062
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24=-0.0026133
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24=-0.042372
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24=-0.01789
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24=0.0094655
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24=8.9992e-13
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25=3.398e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25=-8.5036e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25=0.013426
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25=0.67133
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25=-0.0024994
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25=-0.04234
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25=-0.010738
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25=0.0082498
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26=0.010767
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26=2.2544e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26=-1.9863e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26=-6549.3
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26=-0.0015001
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26=-0.075182
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27=-0.070434
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27=0.013952
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27=4.4861e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27=-1.3022e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27=-4386.9
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27=0.045021
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27=-0.0037673
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28=0.13838
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28=-0.002965
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28=-0.070847
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28=0.012299
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28=5.2415e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28=-1.0387e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28=-3794.7
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29=0.30729
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29=-0.0016815
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29=-0.05513
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29=-0.094949
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29=0.015462
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29=3.6786e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29=-5.2354e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29=-0.039616
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30=0.078393
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30=-0.0015803
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30=-0.063682
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30=0.0016468
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30=0.0092175
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30=5.8119e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30=-5.1885e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30=0.029742
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31=0.89812
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31=-0.0028062
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31=-0.043569
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31=-0.013953
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31=0.010068
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31=1.6699e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31=-9.048e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31=0.010209
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32=0.64105
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32=-0.0024859
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32=-0.042752
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32=-0.011167
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32=0.0083898
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32=4.1984e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32=-8.083e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32=0.014055
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33=-6258.4
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33=0.41317
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33=-0.0018508
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33=-0.076436
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33=0.012698
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33=5.6027e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33=-4.7165e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34=-3814.8
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34=0.081892
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34=-0.0028998
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34=-0.062625
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34=0.012313
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34=4.6553e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34=-9.9558e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35=0.060297
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35=-3.0341e-7
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35=4.8533e-6
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35=0.47691
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35=-0.0047552
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35=-1.5657e-18
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35=-0.018229
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35=0.0085856
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35=1.0526e-10
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36=1.1135e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36=-1.3535e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36=-3.5283e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36=3.8039e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36=1.1343
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36=-0.0019437
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36=-0.049292
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36=0.005575
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37=-0.00033396
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37=1.9217e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37=-2.255e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37=-0.045281
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37=-3.896e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37=-5.6241e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37=0.21652
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37=-0.0019697
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37=-0.061773
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38=-0.057148
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38=0.0033198
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38=3.8609e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38=2.2592e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38=-0.037876
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38=-1.1356e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38=5.7009e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38=0.29918
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38=-0.0010546
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39=0.64659
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39=-0.0018698
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39=-0.040337
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39=0.0049568
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39=3.2087e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39=-9.6364e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39=-1.898e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39=1.3709e-7
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40=-0.034675
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40=-0.0052842
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40=-0.050834
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40=0.0002558
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40=2.2315e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40=-1.8099e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40=-4548.5
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41=-0.0014275
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41=-0.11159
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41=-0.0026503
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41=-3.5998e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41=-5.5996e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41=-517.4
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42=0.03306
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42=-0.0026432
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42=-0.089507
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42=0.004695
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42=1.1034e-10
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42=-5.5006e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42=2232.7
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43=5.1947e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43=3.8406e-7
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43=0.10112
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43=-0.0026021
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43=-0.070766
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43=0.0096967
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43=6.6646e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43=-1.0211e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44=7.5516e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44=2.7039e-7
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44=0.27368
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44=-0.0031423
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44=-0.053714
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44=0.008296
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44=1.98e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44=-1.0118e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45=-4.8683e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45=5.688e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45=0.52552
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45=-0.0018664
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45=-0.051983
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45=0.005428
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45=7.0173e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45=-3.0191e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46=-7.1485e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46=-619.06
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46=-0.28213
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46=-0.0018334
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46=-0.077185
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46=0.0048861
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46=5.6303e-11
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47=5.8354e-11
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47=-8.6209e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47=2826.1
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47=0.083149
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47=-0.0031886
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47=-0.068015
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47=0.011978
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48=0.0054879
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48=-6.0e-10
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48=5.0257e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48=-1780.5
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48=-0.0014629
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48=-0.13041
.include "sky130_fd_pr__pfet_g5v0d10v5.pm3.spice"