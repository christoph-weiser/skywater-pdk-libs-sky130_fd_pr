* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_pfet_01v8_b__toxe_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__overlap_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_b__lint_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__wint_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__rshg_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__xgw_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__dlc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rd_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rs_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_0=0.0073284
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_0=-0.37815
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_0=-0.098732
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_0=0.065703
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_1=-0.0044144
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_1=-0.38258
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_1=0.005625
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_1=-0.016709
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_2=-0.16654
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_2=-0.00075311
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_2=-0.46753
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_2=0.075792
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_3=0.1567
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_3=0.046678
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_3=-0.42184
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_3=-0.42949
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_4=-0.40692
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_4=-0.0027346
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_4=0.0083596
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_4=0.004505
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_5=-0.46458
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_5=0.067987
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_5=-0.14602
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_5=0.00034696
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_6=-0.43843
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_6=-0.90504
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_6=0.18897
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_6=0.05931
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_7=-0.32548
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_7=0.019862
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_7=-0.019001
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_7=0.00046865
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_8=-0.0015768
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_8=-0.37137
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_8=0.0735
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_8=-0.12592
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_0=-0.022271
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_0=-0.34875
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_0=-0.71655
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_0=0.11455
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_0=-0.00043404
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_0=0.025774
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_0=-1656.1
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_1=876.35
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_1=-0.014049
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_1=-0.32181
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_1=0.076806
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_1=-0.008559
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_1=-0.0002533
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_1=0.012035
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_2=-0.0001857
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_2=0.0052953
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_2=15921.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_2=-0.018595
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_2=-0.39574
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_2=1.0073
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_2=-0.1022
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_3=0.12537
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_3=-0.00053503
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_3=0.02819
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_3=-2980.8
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_3=-0.023461
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_3=-0.3112
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_3=-1.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_4=0.011243
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_4=-0.00062465
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_4=0.022876
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_4=-1155.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_4=-0.012789
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_4=-0.32006
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_4=-0.082859
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_5=-0.090506
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_5=0.0077401
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_5=-0.00033445
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_5=9117.5
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_5=-0.018599
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_5=-0.38485
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_5=0.90757
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_6=-0.43115
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_6=-1.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_6=0.15
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_6=0.0058532
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_6=-0.00064602
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_6=-2850.2
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_6=-0.0251
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_7=-0.010953
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_7=-0.29109
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_7=-0.079109
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_7=0.0080531
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_7=0.010416
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_7=-0.00057548
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_7=-3914.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_8=-0.016606
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_8=-0.36184
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_8=0.85881
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_8=-0.081587
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_8=0.011621
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_8=-0.00044041
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_8=11410.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_8=0.0
.include "sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"