* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8__toxe_mult=0.948
.param sky130_fd_pr__nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8__overlap_mult=0.94816
.param sky130_fd_pr__nfet_01v8__lint_diff=1.21275e-8
.param sky130_fd_pr__nfet_01v8__wint_diff=-3.2175e-8
.param sky130_fd_pr__nfet_01v8__dlc_diff=12.773e-9
.param sky130_fd_pr__nfet_01v8__dwc_diff=-3.2175e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_0=-1.1625e-19
.param sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_0=5.3075e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_0=-35091.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_0=0.040393
.param sky130_fd_pr__nfet_01v8__vth0_diff_0=-0.10867
.param sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.99193
.param sky130_fd_pr__nfet_01v8__u0_diff_0=-0.006001
.param sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_1=-5.7353e-20
.param sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_1=3.1406e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_1=-27431.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_1=0.037642
.param sky130_fd_pr__nfet_01v8__vth0_diff_1=-0.078099
.param sky130_fd_pr__nfet_01v8__nfactor_diff_1=1.041
.param sky130_fd_pr__nfet_01v8__u0_diff_1=-0.0051246
.param sky130_fd_pr__nfet_01v8__nfactor_diff_2=1.2221
.param sky130_fd_pr__nfet_01v8__u0_diff_2=0.00091513
.param sky130_fd_pr__nfet_01v8__vth0_diff_2=-0.0069074
.param sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_2=2.7806e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_2=2.1701e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_2=-0.18927
.param sky130_fd_pr__nfet_01v8__a0_diff_2=0.4
.param sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_2=-0.0045103
.param sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_3=-0.0040338
.param sky130_fd_pr__nfet_01v8__nfactor_diff_3=0.90771
.param sky130_fd_pr__nfet_01v8__u0_diff_3=0.00015125
.param sky130_fd_pr__nfet_01v8__vth0_diff_3=-0.013159
.param sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_3=2.5047e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_3=-3.3276e-13
.param sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_3=-0.070457
.param sky130_fd_pr__nfet_01v8__a0_diff_3=0.13825
.param sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_4=0.0042246
.param sky130_fd_pr__nfet_01v8__nfactor_diff_4=1.0788
.param sky130_fd_pr__nfet_01v8__u0_diff_4=-0.0015927
.param sky130_fd_pr__nfet_01v8__vth0_diff_4=-0.015085
.param sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_4=1.1584e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_4=6.7133e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_4=-0.028272
.param sky130_fd_pr__nfet_01v8__a0_diff_4=0.060814
.param sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_5=0.0056805
.param sky130_fd_pr__nfet_01v8__nfactor_diff_5=0.83107
.param sky130_fd_pr__nfet_01v8__u0_diff_5=-0.0016848
.param sky130_fd_pr__nfet_01v8__vth0_diff_5=-0.010908
.param sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_5=1.177e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_5=7.1008e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_5=-0.034049
.param sky130_fd_pr__nfet_01v8__a0_diff_5=0.059073
.param sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_6=0.038669
.param sky130_fd_pr__nfet_01v8__nfactor_diff_6=1.492
.param sky130_fd_pr__nfet_01v8__u0_diff_6=-0.0061621
.param sky130_fd_pr__nfet_01v8__vth0_diff_6=-0.091488
.param sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_6=-1.6835e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_6=4.536e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_6=-36968.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_7=0.021665
.param sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.84742
.param sky130_fd_pr__nfet_01v8__u0_diff_7=-0.0034651
.param sky130_fd_pr__nfet_01v8__vth0_diff_7=-0.067997
.param sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_7=7.5328e-20
.param sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_7=2.1924e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_7=-35764.0
.param sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_8=1.028e-11
.param sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_8=0.0075414
.param sky130_fd_pr__nfet_01v8__nfactor_diff_8=1.5686
.param sky130_fd_pr__nfet_01v8__u0_diff_8=-0.0013777
.param sky130_fd_pr__nfet_01v8__vth0_diff_8=-0.043813
.param sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_8=3.8454e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_8=-37066.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_9=-1.3217e-20
.param sky130_fd_pr__nfet_01v8__vsat_diff_9=-23454.0
.param sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_9=1.0588e-11
.param sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_9=0.0058993
.param sky130_fd_pr__nfet_01v8__nfactor_diff_9=1.5632
.param sky130_fd_pr__nfet_01v8__u0_diff_9=-0.0025729
.param sky130_fd_pr__nfet_01v8__vth0_diff_9=-0.011525
.param sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_10=0.041517
.param sky130_fd_pr__nfet_01v8__ua_diff_10=2.7907e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_10=-7.431e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_10=-31379.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_10=-0.069966
.param sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_10=1.0586
.param sky130_fd_pr__nfet_01v8__u0_diff_10=-0.004511
.param sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_11=0.90844
.param sky130_fd_pr__nfet_01v8__u0_diff_11=-8.1412e-5
.param sky130_fd_pr__nfet_01v8__ags_diff_11=-0.16008
.param sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_11=-0.0012493
.param sky130_fd_pr__nfet_01v8__ua_diff_11=3.3022e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_11=1.3668e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_11=0.025831
.param sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_11=0.0012222
.param sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_12=1.0714
.param sky130_fd_pr__nfet_01v8__u0_diff_12=-0.0028219
.param sky130_fd_pr__nfet_01v8__ags_diff_12=-0.023677
.param sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_12=0.0029922
.param sky130_fd_pr__nfet_01v8__ua_diff_12=1.1894e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_12=-8.5344e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_12=0.03384
.param sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_12=-0.011332
.param sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_13=1.4703
.param sky130_fd_pr__nfet_01v8__u0_diff_13=-0.0040635
.param sky130_fd_pr__nfet_01v8__ags_diff_13=0.011298
.param sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_13=0.0052932
.param sky130_fd_pr__nfet_01v8__ua_diff_13=1.5958e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_13=-1.9512e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_13=0.014103
.param sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_13=-0.014516
.param sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_14=1.1989
.param sky130_fd_pr__nfet_01v8__u0_diff_14=-0.0029321
.param sky130_fd_pr__nfet_01v8__ags_diff_14=-0.0095841
.param sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_14=0.0064914
.param sky130_fd_pr__nfet_01v8__ua_diff_14=1.1147e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_14=-1.3332e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_14=0.035541
.param sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_14=-0.0089431
.param sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_15=-26551.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_15=-0.090092
.param sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_15=1.1928
.param sky130_fd_pr__nfet_01v8__u0_diff_15=-0.0073153
.param sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_15=0.047342
.param sky130_fd_pr__nfet_01v8__ua_diff_15=4.014e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_15=-4.9615e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_16=-24194.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_16=-0.045047
.param sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.54872
.param sky130_fd_pr__nfet_01v8__u0_diff_16=-0.0031346
.param sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_16=0.033945
.param sky130_fd_pr__nfet_01v8__ua_diff_16=1.9692e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_16=4.519e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_17=-23827.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_17=-0.035942
.param sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_17=1.25
.param sky130_fd_pr__nfet_01v8__u0_diff_17=-0.00047656
.param sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_17=0.016135
.param sky130_fd_pr__nfet_01v8__ua_diff_17=3.0188e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_17=1.7684e-19
.param sky130_fd_pr__nfet_01v8__ub_diff_18=1.0996e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_18=-9502.5
.param sky130_fd_pr__nfet_01v8__vth0_diff_18=-0.01712
.param sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_18=0.93684
.param sky130_fd_pr__nfet_01v8__u0_diff_18=-0.0013645
.param sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_18=0.0045237
.param sky130_fd_pr__nfet_01v8__ua_diff_18=6.0012e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_19=1.0534e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_19=1.1911e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_19=0.01338
.param sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_19=0.0027696
.param sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.86302
.param sky130_fd_pr__nfet_01v8__u0_diff_19=-0.00044898
.param sky130_fd_pr__nfet_01v8__ags_diff_19=-0.0031687
.param sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_19=0.004879
.param sky130_fd_pr__nfet_01v8__ua_diff_20=1.7846e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_20=-2.4238e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_20=0.031901
.param sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_20=-0.015969
.param sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_20=1.0179
.param sky130_fd_pr__nfet_01v8__u0_diff_20=-0.0040411
.param sky130_fd_pr__nfet_01v8__ags_diff_20=-0.011538
.param sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_20=0.0029706
.param sky130_fd_pr__nfet_01v8__ags_diff_21=-0.034012
.param sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_21=0.0024091
.param sky130_fd_pr__nfet_01v8__ua_diff_21=1.1125e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_21=-1.5169e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_21=0.050141
.param sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_21=-0.010686
.param sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_21=0.81902
.param sky130_fd_pr__nfet_01v8__u0_diff_21=-0.0026598
.param sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_22=1.1736
.param sky130_fd_pr__nfet_01v8__u0_diff_22=-0.0021258
.param sky130_fd_pr__nfet_01v8__ags_diff_22=0.017294
.param sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_22=0.0068712
.param sky130_fd_pr__nfet_01v8__ua_diff_22=8.0644e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_22=-6.0978e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_22=0.0028956
.param sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_22=-0.0065592
.param sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_23=1.5918
.param sky130_fd_pr__nfet_01v8__u0_diff_23=-0.0025309
.param sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_23=0.038594
.param sky130_fd_pr__nfet_01v8__ua_diff_23=1.3169e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_23=-8.3378e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_23=-19734.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_23=-0.071485
.param sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_24=1.5765
.param sky130_fd_pr__nfet_01v8__u0_diff_24=-0.0098305
.param sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_24=0.031749
.param sky130_fd_pr__nfet_01v8__ua_diff_24=5.3365e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_24=-4.9047e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_24=-18507.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_24=-0.061419
.param sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_25=0.99413
.param sky130_fd_pr__nfet_01v8__u0_diff_25=-0.00035965
.param sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_25=0.014701
.param sky130_fd_pr__nfet_01v8__ua_diff_25=2.2831e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_25=1.9499e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_25=-19710.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_25=-0.017685
.param sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_26=-11407.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_26=-0.013166
.param sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_26=1.1139
.param sky130_fd_pr__nfet_01v8__u0_diff_26=-0.0010353
.param sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_26=0.0022571
.param sky130_fd_pr__nfet_01v8__ua_diff_26=3.58e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_26=3.3057e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_27=0.084507
.param sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_27=-0.013193
.param sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_27=0.95703
.param sky130_fd_pr__nfet_01v8__u0_diff_27=-0.001564
.param sky130_fd_pr__nfet_01v8__ags_diff_27=-0.075834
.param sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_27=0.003712
.param sky130_fd_pr__nfet_01v8__ua_diff_27=7.7409e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_27=3.1147e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_28=0.005117
.param sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_28=-0.0059123
.param sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_28=0.9391
.param sky130_fd_pr__nfet_01v8__u0_diff_28=-0.0015284
.param sky130_fd_pr__nfet_01v8__ags_diff_28=0.0069276
.param sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_28=0.0043703
.param sky130_fd_pr__nfet_01v8__ua_diff_28=6.5911e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_28=1.4716e-20
.param sky130_fd_pr__nfet_01v8__ub_diff_29=5.7406e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_29=-0.031005
.param sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_29=-0.0089838
.param sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.84229
.param sky130_fd_pr__nfet_01v8__u0_diff_29=-0.0011415
.param sky130_fd_pr__nfet_01v8__ags_diff_29=0.030935
.param sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_29=0.0021451
.param sky130_fd_pr__nfet_01v8__ua_diff_29=4.9559e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_30=-2.815e-21
.param sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_30=-0.005506
.param sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_30=9.4355e-5
.param sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.7784
.param sky130_fd_pr__nfet_01v8__u0_diff_30=-0.0010835
.param sky130_fd_pr__nfet_01v8__ags_diff_30=0.018208
.param sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_30=0.0043056
.param sky130_fd_pr__nfet_01v8__ua_diff_30=4.0515e-12
.param sky130_fd_pr__nfet_01v8__ua_diff_31=1.7239e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_31=1.8943e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_31=-14812.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_31=-0.048201
.param sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_31=-0.058235
.param sky130_fd_pr__nfet_01v8__u0_diff_31=0.00031791
.param sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_31=0.032412
.param sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_32=0.030209
.param sky130_fd_pr__nfet_01v8__ua_diff_32=4.6597e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_32=-3.6939e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_32=-17879.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_32=-0.051364
.param sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_32=1.4588
.param sky130_fd_pr__nfet_01v8__u0_diff_32=-0.0082299
.param sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_33=0.69099
.param sky130_fd_pr__nfet_01v8__u0_diff_33=-0.000468
.param sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_33=0.01592
.param sky130_fd_pr__nfet_01v8__ua_diff_33=3.2229e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_33=1.4018e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_33=-20786.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_33=-0.01658
.param sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_34=1.0312
.param sky130_fd_pr__nfet_01v8__u0_diff_34=-0.0010308
.param sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_34=0.0023487
.param sky130_fd_pr__nfet_01v8__ua_diff_34=3.7206e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_34=2.9272e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_34=-8888.2
.param sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_34=-0.015053
.param sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_35=9.7159e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_35=2.515
.param sky130_fd_pr__nfet_01v8__u0_diff_35=-0.003834
.param sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_35=0.0033794
.param sky130_fd_pr__nfet_01v8__ua_diff_35=1.5064e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_35=9.0683e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_35=-0.047761
.param sky130_fd_pr__nfet_01v8__b0_diff_35=1.8786e-8
.param sky130_fd_pr__nfet_01v8__b0_diff_36=9.1484e-8
.param sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_36=1.6098e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_36=0.98042
.param sky130_fd_pr__nfet_01v8__u0_diff_36=-0.002233
.param sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_36=0.0010001
.param sky130_fd_pr__nfet_01v8__ua_diff_36=8.3058e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_36=1.181e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_36=-0.0057401
.param sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_37=-0.066137
.param sky130_fd_pr__nfet_01v8__b0_diff_37=1.8557e-7
.param sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_37=1.5528e-8
.param sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_37=1.8673
.param sky130_fd_pr__nfet_01v8__u0_diff_37=-0.0051091
.param sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_37=0.0048975
.param sky130_fd_pr__nfet_01v8__ua_diff_37=2.335e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_37=-2.9837e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_38=-0.041505
.param sky130_fd_pr__nfet_01v8__b0_diff_38=9.9093e-8
.param sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_38=1.362e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_38=1.4073
.param sky130_fd_pr__nfet_01v8__u0_diff_38=-0.0036085
.param sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_38=0.0098745
.param sky130_fd_pr__nfet_01v8__ua_diff_38=1.4848e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_38=1.0787e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_39=-0.0082635
.param sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_39=1.1142e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_39=1.5277e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_39=0.9461
.param sky130_fd_pr__nfet_01v8__u0_diff_39=-0.0027345
.param sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_39=-0.0017247
.param sky130_fd_pr__nfet_01v8__ua_diff_39=1.0828e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_39=7.0155e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_40=-57437.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_40=-0.14897
.param sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_40=-2.5003e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_40=2.2838e-8
.param sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_40=1.2701
.param sky130_fd_pr__nfet_01v8__u0_diff_40=-0.0010145
.param sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_40=0.033085
.param sky130_fd_pr__nfet_01v8__ua_diff_40=1.9284e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_40=8.61e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_41=2.6772e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_41=-9474.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_41=-0.13141
.param sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_41=1.0704e-6
.param sky130_fd_pr__nfet_01v8__voff_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_41=1.6377e-8
.param sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_41=0.69719
.param sky130_fd_pr__nfet_01v8__u0_diff_41=-0.006133
.param sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_41=0.016032
.param sky130_fd_pr__nfet_01v8__ua_diff_41=4.4403e-11
.param sky130_fd_pr__nfet_01v8__ua_diff_42=1.515e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_42=1.7745e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_42=6287.8
.param sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_42=-0.045618
.param sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_42=3.4771e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_42=5.442e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_42=1.724
.param sky130_fd_pr__nfet_01v8__u0_diff_42=-0.0033408
.param sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_42=0.0094315
.param sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_43=0.011586
.param sky130_fd_pr__nfet_01v8__ua_diff_43=2.0363e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_43=2.8166e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_43=-0.025181
.param sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_43=2.9678e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_43=7.2562e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_43=2.0375
.param sky130_fd_pr__nfet_01v8__u0_diff_43=-0.00084089
.param sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_44=1.5325
.param sky130_fd_pr__nfet_01v8__u0_diff_44=-0.0063868
.param sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_44=0.0039682
.param sky130_fd_pr__nfet_01v8__ua_diff_44=2.7076e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_44=-2.4014e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_44=-0.039391
.param sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_44=2.0206e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_44=5.7041e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_45=1.49
.param sky130_fd_pr__nfet_01v8__u0_diff_45=-0.0039817
.param sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_45=0.0054607
.param sky130_fd_pr__nfet_01v8__ua_diff_45=1.6328e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_45=-3.3128e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_45=-0.022827
.param sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_45=1.4014e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_45=3.2239e-9
.param sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_46=7.6808e-10
.param sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_46=0.64977
.param sky130_fd_pr__nfet_01v8__u0_diff_46=-0.0017403
.param sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_46=0.0020875
.param sky130_fd_pr__nfet_01v8__ua_diff_46=7.7949e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_46=1.8699e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_46=-0.0063547
.param sky130_fd_pr__nfet_01v8__b0_diff_46=9.4853e-8
.param sky130_fd_pr__nfet_01v8__b0_diff_47=4.5808e-7
.param sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_47=1.6807e-8
.param sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_47=1.1215
.param sky130_fd_pr__nfet_01v8__u0_diff_47=-0.0059137
.param sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_47=0.035099
.param sky130_fd_pr__nfet_01v8__ua_diff_47=1.3878e-10
.param sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_47=-1.9739e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_47=-47947.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_47=-0.15378
.param sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_48=-53290.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_48=-0.04144
.param sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_48=1.6886
.param sky130_fd_pr__nfet_01v8__u0_diff_48=-0.00069694
.param sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_48=0.0019981
.param sky130_fd_pr__nfet_01v8__ua_diff_48=6.8934e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_48=2.4766e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_49=-36934.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_49=-0.093996
.param sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.94211
.param sky130_fd_pr__nfet_01v8__u0_diff_49=-0.0040145
.param sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_49=0.03981
.param sky130_fd_pr__nfet_01v8__ua_diff_49=3.2111e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_49=2.0511e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_50=-31469.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_50=-0.12205
.param sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_50=5.7064e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_50=-8.1551e-10
.param sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.571
.param sky130_fd_pr__nfet_01v8__u0_diff_50=-0.0053284
.param sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_50=0.035308
.param sky130_fd_pr__nfet_01v8__ua_diff_50=3.754e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_50=3.2112e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_51=-38324.63321946
.param sky130_fd_pr__nfet_01v8__kt1_diff_51=6.07518e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_51=-0.10491489
.param sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_51=3.22831e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_51=-4.61362e-10
.param sky130_fd_pr__nfet_01v8__voff_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_51=0.00033347
.param sky130_fd_pr__nfet_01v8__u0_diff_51=-0.0019502
.param sky130_fd_pr__nfet_01v8__nfactor_diff_51=0.34959259
.param sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_51=0.03502317
.param sky130_fd_pr__nfet_01v8__ua_diff_51=2.4186e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_51=1.66053e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_51=-4.85723e-17
.param sky130_fd_pr__nfet_01v8__ub_diff_52=4.16095e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_52=3.2537e-5
.param sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_52=-65067.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_52=-0.12224
.param sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_52=-7.39989e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_52=2.7011e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_52=0.00091873
.param sky130_fd_pr__nfet_01v8__u0_diff_52=-0.0083504
.param sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.5935569
.param sky130_fd_pr__nfet_01v8__keta_diff_52=0.00306555
.param sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_52=0.020341
.param sky130_fd_pr__nfet_01v8__ua_diff_52=-4.02468e-11
.param sky130_fd_pr__nfet_01v8__ua_diff_53=-4.99625e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_53=3.05799e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_53=1.15988e-5
.param sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_53=-59191.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_53=-0.12953
.param sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_53=-4.77112e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_53=2.47721e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_53=0.00032751
.param sky130_fd_pr__nfet_01v8__u0_diff_53=-0.0072906
.param sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.56383409
.param sky130_fd_pr__nfet_01v8__keta_diff_53=0.0010928
.param sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_53=0.022274
.param sky130_fd_pr__nfet_01v8__keta_diff_54=-0.00037717
.param sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_54=0.029985
.param sky130_fd_pr__nfet_01v8__ua_diff_54=1.04128e-10
.param sky130_fd_pr__nfet_01v8__ub_diff_54=-6.43431e-20
.param sky130_fd_pr__nfet_01v8__eta0_diff_54=-4.00316e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_54=-49054.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_54=-0.15398
.param sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_54=3.24896e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_54=1.79413e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_54=-0.00011304
.param sky130_fd_pr__nfet_01v8__u0_diff_54=-0.00048232
.param sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.49466752
.param sky130_fd_pr__nfet_01v8__pclm_diff_55=-4.18441e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_55=-0.00096228
.param sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.48878058
.param sky130_fd_pr__nfet_01v8__keta_diff_55=-0.00013962
.param sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_55=0.031175
.param sky130_fd_pr__nfet_01v8__ua_diff_55=1.16564e-10
.param sky130_fd_pr__nfet_01v8__ub_diff_55=-1.09034e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_55=-1.48189e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_55=-47873.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_55=-0.14959
.param sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_55=4.15269e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_55=1.71716e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_56=-7.83128e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_56=0.00065384
.param sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.48174064
.param sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_56=0.030661
.param sky130_fd_pr__nfet_01v8__ua_diff_56=8.51462e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_56=4.16055e-20
.param sky130_fd_pr__nfet_01v8__eta0_diff_56=2.77352e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_56=-48118.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_56=-3.99555e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_56=-0.14576
.param sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_56=2.90133e-7
.param sky130_fd_pr__nfet_01v8__b1_diff_56=1.0645e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_57=6.86799e-9
.param sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_57=-8.11826e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_57=0.001579
.param sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.47867486
.param sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_57=0.030486
.param sky130_fd_pr__nfet_01v8__ua_diff_57=6.22602e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_57=1.46466e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_57=2.87515e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_57=-49294.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_57=-4.14197e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_57=-0.14144
.param sky130_fd_pr__nfet_01v8__b0_diff_57=1.87189e-7
.param sky130_fd_pr__nfet_01v8__b0_diff_58=1.38166e-7
.param sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_58=5.06931e-9
.param sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_58=-7.0636e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_58=0.0016663
.param sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.47711421
.param sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_58=0.03038
.param sky130_fd_pr__nfet_01v8__ua_diff_58=5.13586e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_58=1.96251e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_58=2.50164e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_58=-49772.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_58=-3.60388e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_58=-0.14016
.param sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_59=-42486.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_59=-0.13818
.param sky130_fd_pr__nfet_01v8__b0_diff_59=3.66155e-8
.param sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_59=-5.23278e-11
.param sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_59=8.25295e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_59=0.0016984
.param sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.45856873
.param sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_59=0.0299
.param sky130_fd_pr__nfet_01v8__ua_diff_59=2.10287e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_59=3.16657e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_59=-4.84694e-17
.param sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_60=-41425.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_60=-0.095911
.param sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_60=3.66155e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_60=-5.23278e-11
.param sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_60=8.25291e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_60=0.00078095
.param sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.45856873
.param sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_60=0.012547
.param sky130_fd_pr__nfet_01v8__ua_diff_60=2.10287e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_60=3.16657e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_60=-2.39546e-11
.param sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_61=-37582.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_61=-0.047403
.param sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__u0_diff_61=0.0030431
.param sky130_fd_pr__nfet_01v8__nfactor_diff_61=0.4633
.param sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_61=0.0058357
.param sky130_fd_pr__nfet_01v8__ua_diff_61=-9.108e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_61=4.60449e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_62=-49521.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_62=-0.037598
.param sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_62=5.45502e-17
.param sky130_fd_pr__nfet_01v8__b1_diff_62=-2.18149e-18
.param sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__u0_diff_62=0.0014459
.param sky130_fd_pr__nfet_01v8__nfactor_diff_62=0.0317
.param sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_62=-0.0023861
.param sky130_fd_pr__nfet_01v8__ua_diff_62=2.9602e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_62=2.5142e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8__sf.pm3.spice"