* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param tol_nfom=-0.069u
.param tol_pfom=-0.060u
.param tol_nw=-0.069u
.param tol_poly=-0.041u
.param tol_li=-0.020u
.param tol_m1=-0.025u
.param tol_m2=-0.025u
.param tol_m3=-0.065u
.param tol_m4=-0.065u
.param tol_m5=-0.17u
.param tol_rdl=-1.0u
.param rcn=345
.param rcp=870
.param rdn=132
.param rdp=228
.param rdn_hv=126
.param rdp_hv=222
.param rp1=55.80
.param rnw=2160
.param rl1=14.8
.param rm1=0.145
.param rm2=0.145
.param rm3=0.056
.param rm4=0.056
.param rm5=0.0358
.param rrdl=0.0067
.param rcp1=243.28
.param rcl1=22.6
.param rcvia=15
.param rcvia2=8
.param rcvia3=8
.param rcvia4=0.891
.param rcrdlcon=0.0077
.param rspwres=4829
.param crpf_precision=8.09e-5
.param crpfsw_precision_1_1=4.51e-11
.param crpfsw_precision_2_1=4.86e-11
.param crpfsw_precision_4_1=5.28e-11
.param crpfsw_precision_8_2=5.79e-11
.param crpfsw_precision_16_2=6.36e-11
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/fast.spice"