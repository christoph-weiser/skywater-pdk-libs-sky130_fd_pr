* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__slope=0.0
.subckt sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1 c0 c1 b
.param mult=1.0
.param ctot_a='96.986e-15*sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor+1/sqrt(mult/0.35298)*sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__slope*96.986e-15*sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor'
.param cli2s='7.433e-15*cli2s_vpp'
.param rat_m3=0.1539
.param rat_m2=0.4074
.param rat_m1=0.4025
.param rat_m12li=0.0362
.param cap_m3='rat_m3*ctot_a'
.param cap_m2='rat_m2*ctot_a'
.param cap_m1='rat_m1*ctot_a'
.param cap_m12li='rat_m12li*ctot_a'
.param lm3=5.05
.param wm3=0.30
.param nfm3=34.0
.param nvia2_c0=104.0
.param nvia2_c1=49.0
.param lm2=5.100
.param wm2=0.140
.param nfm2=76.0
.param nvia_c0=124.0
.param nvia_c1=62.0
.param lm1=5.215
.param wm1=0.140
.param nfm1=72.0
.param nmcon=116.0
rm31 c0 z1 r='rm3*lm3/wm3*(1/3)*(1/nfm3)'
ccmvpp11p5x11p7_m3_lishield z1 c1 c='cap_m3'
rvia2_1 c0 d0 r='rcvia2/nvia2_c0'
rvia2_2 c1 d1 r='rcvia2/nvia2_c1'
rm21 d0 a1 r='rm2*lm2/wm2*(1/3)*(1/nfm2)'
cm2 a1 d1 c='cap_m2'
rvia1 d0 e0 r='rcvia/nvia_c0'
rvia2 d1 e1 r='rcvia/nvia_c1'
rm11 e0 b1 r='rm1*lm1/wm1*(1/3)*(1/nfm1)'
cm1 b1 e1 c='cap_m1'
rmcon e0 f0 r='rcl1/nmcon'
rliw f0 g0 r='rl1'
cli2b g0 b c='cli2s'
cm12li e1 g0 c='cap_m12li'
.ends sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1