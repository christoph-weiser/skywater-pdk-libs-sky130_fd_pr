* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult=9.2429e-1
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult=1.0004e+0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult=8.9176e-1
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff=-1.3619e-9
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_0=-0.0019098
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_0=-0.00025989
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_0=-4140.2
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_0=-0.017838
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_1=-0.0088849
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_1=-0.002597
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_1=0.0006887
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_1=-1709.2
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_2=-0.0018947
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_2=-0.012344
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_2=0.00070107
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_2=-3891.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_3=-0.013074
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_3=-0.011262
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_3=-0.0041387
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_3=-6088.7
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_4=-0.008659
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_4=-0.020003
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_4=-0.0021579
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_4=-1519.6
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_5=-0.0014917
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_5=-0.0074298
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_5=-0.0010425
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_5=-415.88
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_6=-0.020457
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_6=-0.010257
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_6=-0.008363
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_6=-5555.5
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_7=-0.0091424
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_7=-0.01706
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_7=-0.0042397
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_7=-790.25
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_8=-0.0013518
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_8=-0.0069456
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_8=-0.0019193
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_8=-105.44
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_0=-0.017526
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_0=-0.0051133
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_0=-0.0060348
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_0=145.4
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_1=-0.0093978
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_1=-0.010042
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_1=-0.0028136
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_1=-1622.4
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_2=-0.0023374
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_2=-0.017756
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_2=-0.0017253
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_2=2328.3
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_3=-0.014282
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_3=-0.0085151
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_3=-0.0046757
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_3=-6719.9
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_4=-0.0069428
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_4=327.64
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_4=-0.0096416
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_4=-0.017088
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_5=-0.019991
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_5=-0.0042474
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_5=9083.2
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_5=-0.0027118
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_6=-0.01916
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_6=-0.013021
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_6=-0.0061579
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_6=-6431.2
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_7=-0.011438
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_7=-0.018674
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_7=-0.0084514
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_7=-2625.5
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_8=-0.0028374
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_8=-0.0065635
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_8=14190.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_8=-0.024019
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_8=0.0
.include "sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"