* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre=0.0
.subckt sky130_fd_pr__nfet_01v8 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__nfet_01v8__model.0 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.52129956+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.026812991 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.58189 eta0=0.08 etab=-0.07 u0=0.03237873 ua=-7.5961167e-10 ub=1.7358267e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.296936 ags=0.436469 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.1 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.52129956+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.026812991 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.58189 eta0=0.08 etab=-0.07 u0=0.03237873 ua=-7.5961167e-10 ub=1.7358267e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.296936 ags=0.436469 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.2 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.216677013e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-2.927416090e-09 wvth0=-3.681462022e-08 pvth0=2.927454790e-13 k1=5.415460247e-01 lk1=-5.410258407e-09 wk1=-6.803836640e-08 pk1=5.410329931e-13 k2=-2.728362245e-02 lk2=3.742405313e-09 wk2=4.706376752e-08 pk2=-3.742454788e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.049993880e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.140741475e-09 wvoff=-2.692155196e-08 pvoff=2.140769775e-13 nfactor=2.586099017e+00 lnfactor=-3.346960113e-08 wnfactor=-4.209072494e-07 pnfactor=3.347004359e-12 eta0=0.08 etab=-0.07 u0=3.236740976e-02 lu0=9.001719900e-11 wu0=1.132038936e-09 pu0=-9.001838903e-15 ua=-7.592259154e-10 lua=-3.067475044e-18 wua=-3.857597462e-17 pua=3.067515596e-22 ub=1.736242864e-18 lub=-3.309285372e-27 wub=-4.161693466e-26 pub=3.309329120e-31 uc=4.876992667e-11 luc=3.753870973e-18 wuc=4.720795745e-17 puc=-3.753920599e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.289894841e+00 la0=5.599046120e-08 wa0=7.041252428e-07 pa0=-5.599120140e-12 ags=4.369120661e-01 lags=-3.523209293e-09 wags=-4.430720065e-08 pags=3.523255870e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=1.950603759e-24 lb1=1.246367018e-30 wb1=1.567407127e-29 pb1=-1.246383495e-34 keta=-8.287889113e-03 lketa=-4.029304676e-09 wketa=-5.067175858e-08 pketa=4.029357943e-13 dwg=0.0 dwb=0.0 pclm=6.801970356e-02 lpclm=-3.316228880e-07 wpclm=-4.170425488e-06 ppclm=3.316272720e-11 pdiblc1=0.39 pdiblc2=3.074732584e-03 lpdiblc2=-1.012977380e-11 wpdiblc2=-1.273900819e-10 ppdiblc2=1.012990772e-15 pdiblcb=-0.025 drout=0.56 pscbe1=7.580453780e+08 lpscbe1=-2.680752404e+01 wpscbe1=-3.371262527e+02 ppscbe1=2.680787844e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.131869363e-01 lkt1=1.247938830e-09 wkt1=1.569383807e-08 pkt1=-1.247955328e-13 kt2=-4.539674530e-02 lkt2=6.632528732e-10 wkt2=8.340940231e-09 pkt2=-6.632616414e-14 at=140000.0 ute=-1.816360220e+00 lute=2.353932011e-08 wute=2.960259503e-07 pute=-2.353963130e-12 ua1=3.613706280e-10 lua1=1.164900625e-16 wua1=1.464956562e-15 pua1=-1.164916025e-20 ub1=-6.204417884e-19 lub1=-1.525028565e-25 wub1=-1.917846515e-24 pub1=1.525048726e-29 uc1=1.691024595e-11 luc1=-8.592269396e-18 wuc1=-1.080547230e-16 puc1=8.592382985e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.3 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.162579434e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.845130344e-08 wvth0=2.110652363e-08 pvth0=6.384801114e-14 k1=5.305679793e-01 lk1=3.797367057e-08 wk1=1.370175511e-07 pk1=-2.693235914e-13 k2=-1.976964001e-02 lk2=-2.595195915e-08 wk2=-8.679876968e-08 pk2=1.547633386e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.379584720e-01 ldsub=8.710549588e-08 wdsub=2.204181943e-06 pdsub=-8.710664742e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.093592126e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.508876654e-08 wvoff=5.581643455e-08 pvoff=-1.128936993e-13 nfactor=2.524931628e+00 lnfactor=2.082566418e-07 wnfactor=1.729922245e-07 pnfactor=9.999843124e-13 eta0=7.415899507e-02 leta0=2.308295641e-08 weta0=5.841082149e-07 peta0=-2.308326157e-12 etab=-6.489376344e-02 letab=-2.017923923e-08 wetab=-5.106304060e-07 petab=2.017950600e-12 u0=3.241892097e-02 lu0=-1.135489536e-10 wu0=1.083486111e-08 pu0=-4.734623749e-14 ua=-7.780901697e-10 lua=7.148181338e-17 wua=1.341701049e-15 pua=-5.147938984e-21 ub=1.738033714e-18 lub=-1.038651141e-26 wub=-7.667795080e-25 pub=3.196689107e-30 uc=5.868885025e-11 luc=-3.544453469e-17 wuc=-3.252598898e-16 puc=1.096556549e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.400419455e+00 la0=-3.807896638e-07 wa0=-1.109326678e-06 pa0=1.567426049e-12 ags=4.443124842e-01 lags=-3.276878091e-08 wags=-1.365734234e-06 pags=5.574447973e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=4.477460477e-24 lb1=-8.739470033e-30 wb1=-3.134814254e-29 pb1=6.118784381e-35 keta=-1.632055236e-02 lketa=2.771482460e-08 wketa=8.771741134e-08 pketa=-1.439617369e-13 dwg=0.0 dwb=0.0 pclm=-6.063528072e-01 lpclm=2.333417024e-06 wpclm=8.545619479e-06 ppclm=-1.708956930e-11 pdiblc1=0.39 pdiblc2=3.180707274e-03 lpdiblc2=-4.289291370e-10 wpdiblc2=-1.239654383e-08 ppdiblc2=4.949922637e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.036964011e+08 lpscbe1=1.879731649e+02 wpscbe1=6.742525055e+02 ppscbe1=-1.316060655e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.113063833e-01 lkt1=-6.183782893e-09 wkt1=3.356221846e-08 pkt1=-1.954092457e-13 kt2=-4.405309717e-02 lkt2=-4.646684630e-09 wkt2=-1.658028237e-08 pkt2=3.215954194e-14 at=1.381587977e+05 lat=7.276212423e-03 wat=1.841226650e-01 pat=-7.276308614e-7 ute=-1.758475983e+00 lute=-2.052122980e-07 wute=-1.608179776e-06 pute=5.171231302e-12 ua1=6.200429155e-10 lua1=-9.057520355e-16 wua1=-5.180235943e-15 pua1=1.461184975e-20 ub1=-9.431076880e-19 lub1=1.122634382e-24 wub1=5.184211542e-24 pub1=-1.281600103e-29 uc1=-6.292278389e-14 luc1=5.848367361e-17 wuc1=1.714481792e-16 puc1=-2.453239098e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.4 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.274191454e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.334034725e-09 wvth0=-1.169960907e-07 pvth0=3.334078801e-13 k1=5.524414795e-01 lk1=-4.720798860e-09 wk1=-2.428261577e-07 pk1=4.720861269e-13 k2=-3.399072719e-02 lk2=1.805910719e-09 wk2=8.501334280e-08 pk2=-1.805934593e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.825849097e-01 wdsub=-2.258520825e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.029702180e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.618209377e-09 wvoff=1.321175511e-07 pvoff=-2.618243989e-13 nfactor=2.623186433e+00 lnfactor=1.647495324e-08 wnfactor=1.529376869e-06 pnfactor=-1.647517103e-12 eta0=8.613056143e-02 leta0=-2.841165134e-10 weta0=-6.130642477e-07 peta0=2.841202694e-14 etab=-7.521863285e-02 letab=-2.632280155e-11 wetab=5.218701842e-07 petab=2.632314954e-15 u0=3.205281457e-02 lu0=6.010471727e-10 wu0=1.737177312e-08 pu0=-6.010551185e-14 ua=-7.785202275e-10 lua=7.232123499e-17 wua=2.409532604e-15 pua=-7.232219108e-21 ub=1.763998182e-18 lub=-6.106606265e-26 wub=-2.257648002e-24 pub=6.106686994e-30 uc=3.956649379e-11 luc=1.880029566e-18 wuc=3.328550213e-16 puc=-1.880054420e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.145470791e+04 lvsat=-2.839416724e-03 wvsat=-1.454727138e-01 pvsat=2.839454261e-7 a0=1.196986241e+00 la0=1.628776154e-08 wa0=5.281828507e-07 pa0=-1.628797687e-12 ags=4.484984837e-01 lags=-4.093935374e-08 wags=-6.072563982e-07 pags=4.093989496e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.775472469e-03 lketa=9.083964511e-09 wketa=4.793635840e-07 pketa=-9.084084601e-13 dwg=0.0 dwb=0.0 pclm=5.771171562e-01 lpclm=2.342448861e-08 wpclm=9.902974737e-07 ppclm=-2.342479828e-12 pdiblc1=4.127280195e-01 lpdiblc1=-4.436238950e-08 wpdiblc1=-2.272832000e-06 ppdiblc1=4.436297597e-12 pdiblc2=2.903550064e-03 lpdiblc2=1.120487551e-10 wpdiblc2=1.870384087e-08 ppdiblc2=-1.120502363e-14 pdiblcb=-2.322221739e-02 lpdiblcb=-3.470020103e-09 wpdiblcb=-1.777806115e-07 ppdiblcb=3.470065977e-13 drout=5.385018536e-01 ldrout=4.196182351e-08 wdrout=2.149843061e-06 pdrout=-4.196237825e-12 pscbe1=7.613803400e+08 lpscbe1=7.538098066e+01 wpscbe1=3.862017059e+03 ppscbe1=-7.538197720e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.170338738e-07 lalpha0=-3.650678645e-13 walpha0=-1.870363463e-11 palpha0=3.650726907e-17 alpha1=8.524364566e-01 lalpha1=-4.755673331e-09 walpha1=-2.436488803e-07 palpha1=4.755736201e-13 beta0=1.405864287e+01 lbeta0=-3.877272492e-07 wbeta0=-1.986454989e-05 pbeta0=3.877323750e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.107990316e-01 lkt1=-7.174073093e-09 wkt1=-4.341025824e-07 pkt1=7.174167934e-13 kt2=-4.499607811e-02 lkt2=-2.806098057e-09 wkt2=-1.438697910e-07 pkt2=2.806135154e-13 at=1.381907748e+05 lat=7.213796952e-03 wat=1.809249139e-01 pat=-7.213892319e-7 ute=-1.804270971e+00 lute=-1.158259318e-07 wute=-4.892967630e-06 pute=1.158274630e-11 ua1=2.791770821e-10 lua1=-2.404224918e-16 wua1=-1.001184057e-14 pua1=2.404256702e-20 ub1=-4.326222229e-19 lub1=1.262275014e-25 wub1=5.085289514e-24 pub1=-1.262291701e-29 uc1=3.129225227e-11 luc1=-2.717896822e-18 wuc1=-9.348456268e-17 puc1=2.717932753e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.5 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.177743821e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.846632285e-09 wvth0=2.014211533e-07 pvth0=3.031255545e-14 k1=5.409461269e-01 lk1=6.221408851e-09 wk1=9.182971227e-07 pk1=-6.331650624e-13 k2=-2.847301392e-02 lk2=-3.446295709e-09 wk2=-3.766155448e-07 pk2=2.588223078e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.833441369e-01 ldsub=-2.862869940e-07 wdsub=-5.221622723e-06 pdsub=2.820520398e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.008867668e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.350117038e-10 wvoff=-5.195676899e-08 pvoff=-8.660755109e-14 nfactor=2.560936479e+00 lnfactor=7.572950242e-08 wnfactor=-4.725996074e-07 pnfactor=2.581262667e-13 eta0=1.962565494e-01 leta0=-1.051109520e-07 weta0=-4.440805742e-06 peta0=3.671966428e-12 etab=-1.427857108e-01 letab=6.428949494e-08 wetab=9.975008253e-07 petab=-4.501114553e-13 u0=3.421955086e-02 lu0=-1.461427936e-09 wu0=-3.817718977e-08 pu0=-7.229509501e-15 ua=-5.462538609e-10 lua=-1.487687063e-16 wua=-5.262435686e-15 pua=7.058174005e-23 ub=1.586329725e-18 lub=1.080531653e-25 wub=5.053581334e-24 pub=-8.527332975e-31 uc=1.249697727e-11 luc=2.764698802e-17 wuc=2.002750928e-16 puc=-6.180512705e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.912535415e+04 lvsat=-6.221491392e-04 wvsat=8.746574143e-02 pvsat=6.221573640e-8 a0=1.284583065e+00 la0=-6.709399097e-08 wa0=-4.554611055e-06 pa0=3.209417259e-12 ags=2.346915626e-01 lags=1.625793921e-07 wags=2.884055336e-06 pags=7.706761918e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.565884743e-03 lketa=-7.597769333e-10 wketa=-7.223979172e-07 pketa=2.355254795e-13 dwg=0.0 dwb=0.0 pclm=6.386699108e-01 lpclm=-3.516640898e-08 wpclm=-2.646241366e-06 ppclm=1.119072399e-12 pdiblc1=3.860471066e-01 lpdiblc1=-1.896533546e-08 wpdiblc1=3.952945608e-07 ppdiblc1=1.896558618e-12 pdiblc2=1.308035497e-03 lpdiblc2=1.630788757e-09 wpdiblc2=2.263590202e-08 ppdiblc2=-1.494787793e-14 pdiblcb=-2.855556522e-02 lpdiblcb=1.606692369e-09 wpdiblcb=3.555612229e-07 ppdiblcb=-1.606713610e-13 drout=5.988291314e-01 ldrout=-1.546256599e-08 wdrout=-3.882964469e-06 pdrout=1.546277040e-12 pscbe1=8.609660156e+08 lpscbe1=-1.941273183e+01 wpscbe1=-6.096682154e+03 ppscbe1=1.941298846e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.211877697e-08 lalpha0=-2.176071273e-13 walpha0=-3.211920158e-12 palpha0=2.176100041e-17 alpha1=8.451270868e-01 lalpha1=2.201976883e-09 walpha1=4.872977606e-07 palpha1=-2.202005994e-13 beta0=1.379882170e+01 lbeta0=-1.404084083e-07 wbeta0=6.117911204e-06 pbeta0=1.404102645e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.100212873e-01 lkt1=-7.914393111e-09 wkt1=2.870581297e-07 pkt1=3.095761367e-14 kt2=-4.858995592e-02 lkt2=6.148459482e-10 wkt2=2.167724799e-07 pkt2=-6.267501009e-14 at=1.694463854e+05 lat=-2.253782494e-02 wat=-6.798199551e-01 pat=9.793745481e-8 ute=-2.097111601e+00 lute=1.629235004e-07 wute=1.189228885e-05 pute=-4.394820425e-12 ua1=-3.446290069e-10 lua1=3.533666721e-16 wua1=2.468880454e-14 pua1=-8.988317748e-21 ub1=-1.033833435e-19 lub1=-1.871687324e-25 wub1=-1.125116664e-23 pub1=2.927445210e-30 uc1=1.779506188e-11 luc1=1.012982226e-17 wuc1=7.068826605e-16 puc1=-4.900610775e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.6 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.274704895e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.465145582e-09 wvth0=5.927388908e-07 pvth0=-1.465164951e-13 k1=5.714933154e-01 lk1=-7.582285245e-09 wk1=-2.160840107e-06 pk1=7.582385482e-13 k2=-4.035228131e-02 lk2=1.921719520e-09 wk2=6.214277462e-07 pk2=-1.921744925e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.596735873e-01 ldsub=-4.462122378e-09 wdsub=3.264169827e-08 pdsub=4.462181368e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.997113297e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.212541797e-10 wvoff=-1.946532767e-07 pvoff=-2.212571047e-14 nfactor=2.717398776e+00 lnfactor=5.027162994e-09 wnfactor=1.211138394e-06 pnfactor=-5.027229453e-13 eta0=-3.635104429e-02 weta0=3.685153146e-6 etab=-5.499564097e-04 letab=1.586000423e-11 wetab=4.926599094e-09 petab=-1.586021390e-15 u0=3.069161679e-02 lu0=1.327784406e-10 wu0=-2.479200630e-08 pu0=-1.327801959e-14 ua=-9.074470998e-10 lua=1.444765570e-17 wua=-1.908972253e-15 pua=-1.444784669e-21 ub=1.847120339e-18 lub=-9.793157896e-27 wub=9.992793527e-25 pub=9.793287361e-31 uc=7.379078568e-11 luc=-5.051941959e-20 wuc=5.232212330e-17 puc=5.052008746e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.861525495e+04 lvsat=-3.916450013e-04 wvsat=1.384763361e-01 pvsat=3.916501788e-8 a0=1.136105942e+00 wa0=2.547739473e-6 ags=5.196714811e-01 lags=3.380238157e-08 wags=1.207001145e-05 pags=-3.380282844e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.172846096e-03 lketa=3.215917632e-10 wketa=-1.300183284e-07 pketa=-3.215960147e-14 dwg=0.0 dwb=0.0 pclm=5.532722347e-01 lpclm=3.423178290e-09 wpclm=5.877843031e-07 ppclm=-3.423223544e-13 pdiblc1=2.904675970e-01 lpdiblc1=2.422522894e-08 wpdiblc1=9.953371882e-06 ppdiblc1=-2.422554920e-12 pdiblc2=4.863094537e-03 lpdiblc2=2.432512251e-11 wpdiblc2=-5.060180628e-09 ppdiblc2=-2.432544409e-15 pdiblcb=-3.715857107e-02 lpdiblcb=5.494227253e-09 wpdiblcb=1.215873180e-06 ppdiblcb=-5.494299887e-13 drout=5.950831792e-01 ldrout=-1.376984140e-08 wdrout=-3.508364304e-06 pdrout=1.377002343e-12 pscbe1=8.325466090e+08 lpscbe1=-6.570541976e+00 wpscbe1=-3.254703929e+03 ppscbe1=6.570628839e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.237036965e-07 lalpha0=9.230301785e-14 walpha0=6.537123385e-11 palpha0=-9.230423809e-18 alpha1=0.85 beta0=1.350798108e+01 lbeta0=-8.983061558e-09 wbeta0=3.520235693e-05 pbeta0=8.983180315e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.284421631e-01 lkt1=4.096506828e-10 wkt1=4.462222094e-07 pkt1=-4.096560984e-14 kt2=-4.746478522e-02 lkt2=1.064026884e-10 wkt2=1.016213658e-07 pkt2=-1.064040951e-14 at=1.178987885e+05 lat=7.555546764e-04 wat=-2.958827653e-01 pat=-7.555646648e-8 ute=-1.702631217e+00 lute=-1.533469017e-08 wute=-1.226894547e-06 pute=1.533489290e-12 ua1=4.578996562e-10 lua1=-9.280782745e-18 wua1=2.744070655e-15 pua1=9.280905437e-22 ub1=-4.913213252e-19 lub1=-1.186692925e-26 wub1=-7.398965290e-24 pub1=1.186708613e-30 uc1=4.652153009e-11 luc1=-2.851122920e-18 wuc1=-1.008562642e-15 puc1=2.851160611e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.7 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.232755496e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.312024229e-09 wvth0=1.012238420e-06 pvth0=-2.312054794e-13 k1=5.516607773e-01 lk1=-3.578472617e-09 wk1=-1.775600772e-07 pk1=3.578519925e-13 k2=-3.407796028e-02 lk2=6.550533163e-10 wk2=-6.012651373e-09 pk2=-6.550619761e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.150206873e-01 ldsub=4.552449726e-09 wdsub=4.497990729e-06 pdsub=-4.552509909e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.006521549e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.587395722e-10 wvoff=-1.265501813e-07 pvoff=-3.587443148e-14 nfactor=2.818718930e+00 lnfactor=-1.542745090e-08 wnfactor=-8.921010896e-06 pnfactor=1.542765486e-12 eta0=-1.014554357e-01 leta0=1.314333965e-08 weta0=1.019567836e-05 peta0=-1.314351340e-12 etab=-4.367255160e-03 letab=7.865000933e-10 wetab=3.866615206e-07 petab=-7.865104908e-14 u0=3.263354498e-02 lu0=-2.592599658e-10 wu0=-2.189873933e-07 pu0=2.592633933e-14 ua=-6.356208837e-10 lua=-4.042889264e-17 wua=-2.909195322e-14 pua=4.042942711e-21 ub=1.640513751e-18 lub=3.191678652e-26 wub=2.166021120e-23 pub=-3.191720846e-30 uc=7.379740406e-11 luc=-5.185554374e-20 wuc=5.166027706e-17 puc=5.185622927e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.804496936e+04 lvsat=-2.765151772e-04 wvsat=1.955056484e-01 pvsat=2.765188327e-8 a0=1.136105942e+00 wa0=2.547739473e-6 ags=8.616313619e-01 lags=-3.523282112e-08 wags=-2.212642870e-05 pags=3.523328690e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.668458393e-03 lketa=1.965605718e-11 wketa=-2.795815353e-07 pketa=-1.965631703e-15 dwg=0.0 dwb=0.0 pclm=5.524199353e-01 lpclm=3.595241343e-09 wpclm=6.730153688e-07 ppclm=-3.595288872e-13 pdiblc1=4.468764739e-01 lpdiblc1=-7.350751536e-09 wpdiblc1=-5.687722581e-06 ppdiblc1=7.350848712e-13 pdiblc2=5.875679373e-03 lpdiblc2=-1.800965168e-10 wpdiblc2=-1.063200029e-07 ppdiblc2=1.800988977e-14 pdiblcb=9.721065548e-03 lpdiblcb=-3.969880667e-09 wpdiblcb=-3.472152456e-06 ppdiblcb=3.969933149e-13 drout=4.867223816e-01 ldrout=8.106144785e-09 wdrout=7.327858709e-06 pdrout=-8.106251948e-13 pscbe1=7.994179815e+08 lpscbe1=1.174984772e-01 wpscbe1=5.820261965e+01 ppscbe1=-1.175000306e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.395410281e-07 lalpha0=7.531217418e-14 walpha0=5.695485574e-11 palpha0=-7.531316981e-18 alpha1=8.983796825e-01 lalpha1=-9.766938691e-09 walpha1=-4.838032212e-06 palpha1=9.767067810e-13 beta0=1.287813408e+01 lbeta0=1.181710817e-07 wbeta0=9.818789013e-05 pbeta0=-1.181726440e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.217986276e-01 lkt1=-9.315529168e-10 wkt1=-2.181401280e-07 pkt1=9.315652319e-14 kt2=-4.640015474e-02 lkt2=-1.085259792e-10 wkt2=-4.843090487e-09 pkt2=1.085274139e-14 at=1.230656651e+05 lat=-2.875395341e-04 wat=-8.125772537e-01 pat=2.875433354e-8 ute=-1.914121832e+00 lute=2.736124665e-08 wute=1.992244653e-05 pute=-2.736160837e-12 ua1=1.260674364e-10 lua1=5.770983763e-17 wua1=3.592773132e-14 pua1=-5.771060055e-21 ub1=-3.112059696e-19 lub1=-4.822879736e-26 wub1=-2.541073897e-23 pub1=4.822943495e-30 uc1=3.829448063e-11 luc1=-1.190237948e-18 wuc1=-1.858468196e-16 puc1=1.190253682e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.8 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.283993306e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.636294877e-09 wvth0=4.998535529e-07 pvth0=-1.636316508e-13 k1=5.286178406e-01 lk1=-5.395470780e-10 wk1=2.126764059e-06 pk1=5.395542108e-14 k2=-2.743879665e-02 lk2=-2.205262220e-10 wk2=-6.699377910e-07 pk2=2.205291373e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.310270715e-01 ldsub=2.441511775e-09 wdsub=2.897331152e-06 pdsub=-2.441544052e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=4.019416492e-03 lcdscd=1.820727866e-10 wcdscd=1.380602161e-07 pcdscd=-1.820751936e-14 cit=0.0 voff='-1.140387909e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.124182510e-09 wvoff=1.212131113e-06 pvoff=-2.124210592e-13 nfactor=2.386040208e+00 lnfactor=4.163465155e-08 wnfactor=3.434743324e-05 pnfactor=-4.163520196e-12 eta0=-9.516126367e-03 leta0=1.018291590e-09 weta0=1.001625878e-06 peta0=-1.018305051e-13 etab=-2.041762496e-03 letab=4.798117953e-10 wetab=1.541091799e-07 petab=-4.798181384e-14 u0=2.764047574e-02 lu0=3.992309992e-10 wu0=2.803261320e-07 pu0=-3.992362770e-14 ua=-1.369294987e-09 lua=5.632878184e-17 wua=4.427642707e-14 pua=-5.632952651e-21 ub=2.243412957e-18 lub=-4.759416359e-26 wub=-3.863050637e-23 pub=4.759479278e-30 uc=6.489801803e-11 luc=1.121804386e-18 wuc=9.416106454e-16 puc=-1.121819216e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.935779813e+04 lvsat=-4.496523485e-04 wvsat=6.422103564e-02 pvsat=4.496582929e-8 a0=1.136105942e+00 wa0=2.547739473e-6 ags=5.944752050e-01 wags=4.589540168e-6 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.860473495e-02 lketa=-2.082036032e-09 wketa=-1.873230259e-06 pketa=2.082063556e-13 dwg=0.0 dwb=0.0 pclm=5.497838770e-01 lpclm=3.942887345e-09 wpclm=9.366246818e-07 ppclm=-3.942939470e-13 pdiblc1=3.941646009e-01 lpdiblc1=-3.990570185e-10 wpdiblc1=-4.164656001e-07 ppdiblc1=3.990622940e-14 pdiblc2=4.694771318e-03 lpdiblc2=-2.435718152e-11 wpdiblc2=1.177236384e-08 ppdiblc2=2.435750352e-15 pdiblcb=1.694746582e-03 lpdiblcb=-2.911361695e-09 wpdiblcb=-2.669509949e-06 ppdiblcb=2.911400184e-13 drout=5.020872680e-01 ldrout=6.079808207e-09 wdrout=5.791349761e-06 pdrout=-6.079888582e-13 pscbe1=7.989383347e+08 lpscbe1=1.807547819e-01 wpscbe1=1.061679376e+02 ppscbe1=-1.807571715e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.668446184e-08 lalpha0=-6.810196562e-16 walpha0=-6.684550204e-13 palpha0=6.810286593e-20 alpha1=7.371140741e-01 lalpha1=1.150093102e-08 walpha1=1.128874183e-05 palpha1=-1.150108306e-12 beta0=1.348272074e+01 lbeta0=3.843758828e-08 wbeta0=3.772842476e-05 pbeta0=-3.843809643e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.176875281e-01 lkt1=-1.473728829e-09 wkt1=-6.292555120e-07 pkt1=1.473748312e-13 kt2=-4.550306418e-02 lkt2=-2.268351789e-10 wkt2=-9.455333206e-08 pkt2=2.268381776e-14 at=1.200576762e+05 lat=1.091570525e-04 wat=-5.117743852e-01 pat=-1.091584956e-8 ute=-1.240206601e+00 lute=-6.151536793e-08 wute=-4.746996749e-05 pute=6.151618116e-12 ua1=1.213291357e-09 lua1=-8.567434029e-17 wua1=-7.279609809e-14 pua1=8.567547291e-21 ub1=-1.049198629e-18 lub1=4.909841254e-26 wub1=4.838950259e-23 pub1=-4.909906162e-30 uc1=3.621795341e-11 luc1=-9.163834616e-19 wuc1=2.180864725e-17 puc1=9.163955762e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.9 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.189603568e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.338077633e-07 wvth0=1.637751506e-08 pvth0=-1.636963437e-12 k1=5.418246413e-01 lk1=-9.585297950e-08 wk1=-6.714206551e-09 pk1=6.710975742e-13 k2=-2.606591356e-02 lk2=-7.467179492e-08 wk2=-5.230529684e-09 pk2=5.228012806e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.045276656e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.405778430e-08 wvoff=-5.187520128e-09 pvoff=5.185023945e-13 nfactor=2.767435424e+00 lnfactor=-1.854561413e-05 wnfactor=-1.299063258e-06 pnfactor=1.298438162e-10 eta0=0.08 etab=-0.07 u0=3.182751958e-02 lu0=5.509451828e-08 wu0=3.859201639e-09 pu0=-3.857344629e-13 ua=-7.361897331e-10 lua=-2.341066649e-15 wua=-1.639845220e-16 pua=1.639056143e-20 ub=1.668772713e-18 lub=6.702172130e-24 wub=4.694665544e-25 pub=-4.692406518e-29 uc=4.770841727e-11 luc=1.532844783e-16 wuc=1.073710649e-17 puc=-1.073193990e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.318204716e+00 la0=-2.125848135e-06 wa0=-1.489091267e-07 pa0=1.488374731e-11 ags=4.296636097e-01 lags=6.802115605e-07 wags=4.764672876e-08 pags=-4.762380163e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=7.930748498e-25 lb1=1.313635138e-28 wb1=9.201610313e-30 pb1=-9.197182590e-34 keta=-7.168310544e-03 lketa=-1.625506902e-07 wketa=-1.138617615e-08 pketa=1.138069723e-12 dwg=0.0 dwb=0.0 pclm=5.785204888e-02 lpclm=-3.152087405e-06 wpclm=-2.207940329e-07 ppclm=2.206877890e-11 pdiblc1=0.39 pdiblc2=3.148441603e-03 lpdiblc2=-7.494682181e-09 wpdiblc2=-5.249794472e-10 ppdiblc2=5.247268324e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.171647721e+08 lpscbe1=3.749133877e+03 wpscbe1=2.626153028e+02 ppscbe1=-2.624889349e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.201210271e-01 lkt1=7.087614958e-07 wkt1=4.964656397e-08 pkt1=-4.962267454e-12 kt2=-4.543567811e-02 lkt2=1.222822406e-08 wkt2=8.565495046e-10 pkt2=-8.561373415e-14 at=140000.0 ute=-1.857243378e+00 lute=4.382228070e-06 wute=3.069616048e-07 pute=-3.068138980e-11 ua1=3.031015403e-10 lua1=7.288337211e-15 wua1=5.105256164e-16 pua1=-5.102799566e-20 ub1=-5.512035611e-19 lub1=-8.837389381e-24 wub1=-6.190319590e-25 pub1=6.187340870e-29 uc1=1.657636884e-11 luc1=-7.462965572e-17 wuc1=-5.227577962e-18 puc1=5.225062504e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.10 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.306789393e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=-6.566805431e-8 k1=5.370204336e-01 wk1=2.692159822e-8 k2=-2.980850781e-02 wk2=2.097257771e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.082394853e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=2.080012457e-8 nfactor=1.837918346e+00 wnfactor=5.208785109e-6 eta0=0.08 etab=-0.07 u0=3.458888921e-02 wu0=-1.547403631e-8 ua=-8.535253692e-10 wua=6.575200484e-16 ub=2.004689519e-18 wub=-1.882395166e-24 uc=5.539112540e-11 wuc=-4.305200694e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.211655958e+00 wa0=5.970730348e-7 ags=4.637562128e-01 wags=-1.910465635e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=7.377091353e-24 wb1=-3.689520928e-29 keta=-1.531544666e-02 wketa=4.565454715e-8 dwg=0.0 dwb=0.0 pclm=-1.001324241e-01 wpclm=8.853061337e-7 pdiblc1=0.39 pdiblc2=2.772803728e-03 wpdiblc2=2.104982271e-9 pdiblcb=-0.025 drout=0.56 pscbe1=9.050735651e+08 wpscbe1=-1.052994664e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.845974844e-01 wkt1=-1.990651968e-7 kt2=-4.482279233e-02 wkt2=-3.434461160e-9 at=140000.0 ute=-1.637603532e+00 wute=-1.230807681e-6 ua1=6.683972841e-10 wua1=-2.047027512e-15 ub1=-9.941387100e-19 wub1=2.482099644e-24 uc1=1.283588664e-11 wuc1=2.096074235e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.11 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.352278362e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.617228753e-08 wvth0=-1.317534910e-07 pvth0=5.255035288e-13 k1=5.247225531e-01 lk1=9.779128238e-08 wk1=4.974817533e-08 pk1=-1.815142248e-13 k2=-2.539121550e-02 lk2=-3.512578278e-08 wk2=3.381441707e-08 pk2=-1.021167784e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.176657393e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.495645024e-08 wvoff=6.175965188e-08 pvoff=-3.257052870e-13 nfactor=1.003826239e+00 lnfactor=6.632601178e-06 wnfactor=1.065709396e-05 pnfactor=-4.332430364e-11 eta0=0.08 etab=-0.07 u0=3.655933359e-02 lu0=-1.566873923e-08 wu0=-2.821696961e-08 pu0=1.013302892e-13 ua=-8.955188119e-10 lua=3.339268589e-16 wua=9.156544803e-16 pua=-2.052654284e-21 ub=2.189901814e-18 lub=-1.472786132e-24 wub=-3.217829322e-24 pub=1.061921349e-29 uc=1.758025073e-10 luc=-9.574969798e-16 wuc=-8.421880439e-16 puc=6.354634669e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.567580345e+00 la0=-2.830268373e-06 wa0=-1.240040390e-06 pa0=1.460850734e-11 ags=6.188908391e-01 lags=-1.233612087e-06 wags=-1.318399187e-06 pags=8.964573908e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=1.466543814e-23 lb1=-5.795606635e-29 wb1=-7.334657842e-29 pb1=2.898569497e-34 keta=-2.853553507e-02 lketa=1.051245699e-07 wketa=9.108853054e-08 pketa=-3.612856292e-13 dwg=0.0 dwb=0.0 pclm=-1.018047063e+00 lpclm=7.299147977e-06 wpclm=3.433477658e-06 ppclm=-2.026275673e-11 pdiblc1=0.39 pdiblc2=2.812183000e-03 lpdiblc2=-3.131392862e-10 wpdiblc2=1.710804096e-09 ppdiblc2=3.134457937e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.006242765e+09 lpscbe1=-8.044854355e+02 wpscbe1=-2.074836076e+03 ppscbe1=8.125561314e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.593635450e-01 lkt1=-2.006572832e-07 wkt1=-3.611410554e-07 pkt1=1.288807940e-12 kt2=-3.211876938e-02 lkt2=-1.010208787e-07 wkt2=-8.462244468e-08 pkt2=6.455971836e-13 at=140000.0 ute=-1.116766532e+00 lute=-4.141633839e-06 wute=-4.602054729e-06 pute=2.680775535e-11 ua1=1.924027327e-09 lua1=-9.984620684e-15 wua1=-9.475706166e-15 pua1=5.907196864e-20 ub1=-2.197589049e-18 lub1=9.569693889e-24 wub1=9.124269302e-24 pub1=-5.281774270e-29 uc1=-2.775741172e-11 luc1=3.227930779e-16 wuc1=2.046779313e-16 puc1=-1.460897224e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.12 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.127732553e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.256554436e-08 wvth0=4.550394741e-08 pvth0=-1.749967743e-13 k1=5.754419082e-01 lk1=-1.026455734e-07 wk1=-1.771592746e-07 pk1=7.151970154e-13 k2=-4.465406786e-02 lk2=4.099871750e-08 wk2=8.742512252e-08 pk2=-3.139799067e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.873006811e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.939387901e-08 wvoff=-8.861484891e-08 pvoff=2.685568456e-13 nfactor=2.787565788e+00 lnfactor=-4.165252560e-07 wnfactor=-1.665794101e-06 pnfactor=5.374283558e-12 eta0=1.575872698e-01 leta0=-3.066156572e-7 etab=-1.378255040e-01 letab=2.680383207e-07 wetab=-1.180622676e-11 petab=4.665680321e-17 u0=3.464830930e-02 lu0=-8.116598640e-09 wu0=-4.773804483e-09 pu0=8.685690340e-15 ua=-4.140529290e-10 lua=-1.568769016e-15 wua=-1.207040894e-15 pua=6.335985233e-21 ub=1.384924306e-18 lub=1.708389185e-24 wub=1.705453154e-24 pub=-8.837012986e-30 uc=-2.099467880e-10 luc=5.669383311e-16 wuc=1.555544714e-15 puc=-3.120919862e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=5.419979687e-01 la0=1.222711135e-06 wa0=4.900758562e-06 pa0=-9.659199367e-12 ags=-8.205227586e-02 lags=1.536431691e-06 wags=2.319514941e-06 pags=-5.412029814e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.736793793e-06 lketa=-7.625749729e-09 wketa=-2.651486715e-08 pketa=1.034690036e-13 dwg=0.0 dwb=0.0 pclm=8.366832526e-01 lpclm=-3.052551792e-08 wpclm=-1.557540633e-06 ppclm=-5.388463726e-13 pdiblc1=0.39 pdiblc2=1.346592463e-03 lpdiblc2=5.478700110e-09 wpdiblc2=4.446845419e-10 ppdiblc2=8.138011748e-15 pdiblcb=-0.025 drout=0.56 pscbe1=8.052807137e+08 lpscbe1=-1.030732470e+01 wpscbe1=-3.697197686e+01 ppscbe1=7.216489917e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.047328192e-01 lkt1=-2.136331085e-08 wkt1=-1.246142074e-08 pkt1=-8.913248269e-14 kt2=-5.824718564e-02 lkt2=2.235513037e-09 wkt2=8.279710150e-08 pkt2=-1.602493999e-14 at=1.674588794e+05 lat=-1.085142239e-01 wat=-2.101664194e-02 pat=8.305526796e-8 ute=-2.534042581e+00 lute=1.459272449e-06 wute=3.821811709e-06 pute=-6.482362377e-12 ua1=-1.722122763e-09 lua1=4.424530583e-15 wua1=1.121802015e-14 pua1=-2.270717521e-20 ub1=1.240325910e-18 lub1=-4.016536919e-24 wub1=-1.010271014e-23 pub1=2.316499205e-29 uc1=6.749233604e-11 luc1=-5.362259045e-17 wuc1=-3.015279406e-16 puc1=5.395681432e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.13 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.278145439e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.320673879e-08 wvth0=-1.197644029e-07 pvth0=1.475873786e-13 k1=4.355608814e-01 lk1=1.703855450e-07 wk1=5.754925450e-07 pk1=-7.538897709e-13 k2=1.065032698e-02 lk2=-6.694888002e-08 wk2=-2.275330519e-07 pk2=3.007809697e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.119150256e+00 ldsub=-1.676959062e-06 wdsub=-6.015187592e-06 pdsub=1.174093037e-11 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.043752606e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.856325128e-09 wvoff=1.419547061e-07 pvoff=-1.814874881e-13 nfactor=2.353536152e+00 lnfactor=4.306489445e-07 wnfactor=3.417285318e-06 pnfactor=-4.547282580e-12 eta0=-6.282989008e-03 leta0=1.323958737e-08 weta0=3.395277610e-08 peta0=-6.627177857e-14 etab=-9.542264724e-04 letab=8.818745641e-10 wetab=1.921162046e-09 petab=-3.726267242e-15 u0=3.466541312e-02 lu0=-8.149983252e-09 wu0=-9.198705826e-10 pu0=1.163269984e-15 ua=-9.456722347e-10 lua=-5.311113938e-16 wua=3.579817630e-15 pua=-3.007392968e-21 ub=2.163821122e-18 lub=1.880752899e-25 wub=-5.056937149e-24 pub=4.362368161e-30 uc=7.464307000e-11 luc=1.145279441e-17 wuc=8.727261657e-17 puc=-2.550274511e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.156320532e+04 lvsat=1.140616692e-01 wvsat=2.738469809e-01 pvsat=-5.345167189e-7 a0=2.146402396e+00 la0=-1.908895384e-06 wa0=-6.118985362e-06 pa0=1.185002942e-11 ags=1.388185770e+00 lags=-1.333298016e-06 wags=-7.186309668e-06 pags=1.314220863e-11 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.996480180e-02 lketa=-1.051603427e-07 wketa=8.210665349e-08 pketa=-1.085472787e-13 dwg=0.0 dwb=0.0 pclm=1.093259657e+00 lpclm=-5.313321258e-07 wpclm=-2.623382369e-06 ppclm=1.541549861e-12 pdiblc1=-1.764509983e-01 lpdiblc1=1.105644941e-06 wpdiblc1=1.852200019e-06 ppdiblc1=-3.615274026e-12 pdiblc2=6.759685497e-03 lpdiblc2=-5.087013333e-09 wpdiblc2=-8.294204968e-09 ppdiblc2=2.519528414e-14 pdiblcb=-4.838917727e-02 lpdiblcb=4.565289072e-08 wpdiblcb=-1.578621569e-09 ppdiblcb=3.081281447e-15 drout=8.455643000e-01 ldrout=-5.573875314e-7 pscbe1=2.297844770e+09 lpscbe1=-2.923614748e+03 wpscbe1=-6.895265160e+03 ppscbe1=1.345873706e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=4.019886220e-07 lalpha0=-7.260775235e-13 walpha0=-1.999856238e-11 palpha0=3.903481394e-17 alpha1=8.176360460e-01 lalpha1=6.317058690e-8 beta0=1.188073775e+01 lbeta0=3.863284386e-06 wbeta0=-4.616334817e-06 pbeta0=9.010536218e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.587235025e-01 lkt1=8.402007807e-08 wkt1=-9.856792995e-08 pkt1=7.893717662e-14 kt2=-8.643118763e-02 lkt2=5.724733103e-08 wkt2=1.462307529e-07 pkt2=-1.398398789e-13 at=1.550323615e+05 lat=-8.425913961e-02 wat=6.301154250e-02 pat=-8.095774871e-8 ute=-2.543043770e+00 lute=1.476841699e-06 wute=2.794186225e-07 pute=4.319673833e-13 ua1=-8.183641789e-10 lua1=2.660501373e-15 wua1=-2.327600791e-15 pua1=3.732264941e-21 ub1=-3.640067860e-19 lub1=-8.850704119e-25 wub1=4.604890746e-24 pub1=-5.542494679e-30 uc1=1.242641734e-11 luc1=5.385952999e-17 wuc1=3.860122244e-17 puc1=-1.243235078e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.14 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.488223603e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.209797531e-09 wvth0=-1.595573989e-08 pvth0=4.877388462e-14 k1=7.125364581e-01 lk1=-9.326224387e-08 wk1=-2.830620379e-07 pk1=6.335202399e-14 k2=-1.032796931e-01 lk2=4.149894140e-08 wk2=1.471301038e-07 pk2=-5.585376953e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.668727950e+00 ldsub=9.767692334e-07 wdsub=1.264625573e-05 pdsub=-6.022542955e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.073809901e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.995228284e-09 wvoff=-6.488620375e-09 pvoff=-4.018710599e-14 nfactor=2.743189981e+00 lnfactor=5.974486819e-08 wnfactor=-1.748615061e-06 pnfactor=3.700398380e-13 eta0=-4.283255210e-01 leta0=4.149738547e-07 weta0=-6.790555220e-08 peta0=3.068522884e-14 etab=2.295546556e-04 letab=-2.449441998e-10 wetab=-3.795099185e-09 petab=1.714933215e-15 u0=2.966764624e-02 lu0=-3.392703923e-09 wu0=-6.307839848e-09 pu0=6.291975557e-15 ua=-1.289451303e-09 lua=-2.038746302e-16 wua=-5.907108195e-17 pua=4.563960574e-22 ub=2.327244664e-18 lub=3.251552522e-26 wub=-1.338027262e-25 pub=-3.238699564e-31 uc=8.747918441e-11 luc=-7.656590146e-19 wuc=-3.246994837e-16 puc=1.371209637e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.860802746e+05 lvsat=-4.253900322e-02 wvsat=-6.613600964e-01 pvsat=3.556891290e-7 a0=-1.087194449e+00 la0=1.169104015e-06 wa0=1.205096704e-05 pa0=-5.445603036e-12 ags=-1.153523214e+00 lags=1.086106473e-06 wags=1.260339399e-05 pags=-5.695234280e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-7.987772330e-02 lketa=1.843428994e-08 wketa=-1.381823485e-07 pketa=1.011416368e-13 dwg=0.0 dwb=0.0 pclm=2.789131805e-01 lpclm=2.438288122e-07 wpclm=-1.274686556e-07 ppclm=-8.342629811e-13 pdiblc1=6.969870319e-01 lpdiblc1=2.742358753e-07 wpdiblc1=-1.781695979e-06 ppdiblc1=-1.562374696e-13 pdiblc2=-1.357929454e-03 lpdiblc2=2.639990103e-09 wpdiblc2=4.130118108e-08 ppdiblc2=-2.201362152e-14 pdiblcb=2.177835454e-02 lpdiblcb=-2.113824963e-08 wpdiblcb=3.157243138e-09 ppdiblcb=-1.426698187e-15 drout=9.900807710e-01 ldrout=-6.949500144e-07 wdrout=-6.622243181e-06 pdrout=6.303587461e-12 pscbe1=-1.438980881e+09 lpscbe1=6.333985896e+02 wpscbe1=1.000598665e+04 ppscbe1=-2.629243420e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.960165063e-05 lalpha0=1.831500661e-11 walpha0=1.344604612e-10 palpha0=-1.079917959e-16 alpha1=9.147279080e-01 lalpha1=-2.924931179e-8 beta0=2.189528436e+00 lbeta0=1.308816240e-05 wbeta0=8.739831152e-05 pbeta0=-7.857645735e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.687456453e-01 lkt1=-1.628134625e-09 wkt1=-1.925930815e-09 pkt1=-1.305450616e-14 kt2=-1.802414066e-02 lkt2=-7.868037253e-09 wkt2=2.771365030e-09 pkt2=-3.283613306e-15 at=7.927578925e+04 lat=-1.214789789e-02 wat=-4.850657651e-02 pat=2.519422994e-8 ute=-6.988367146e-01 lute=-2.786239574e-07 wute=2.102516130e-06 pute=-1.303404495e-12 ua1=2.545780189e-09 lua1=-5.417637325e-16 wua1=4.452119043e-15 pua1=-2.721221554e-21 ub1=-1.238079919e-18 lub1=-5.305680410e-26 wub1=-3.306790541e-24 pub1=1.988484417e-30 uc1=1.459532890e-10 luc1=-7.324216211e-17 wuc1=-1.903943543e-16 puc1=9.365303081e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.15 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.899946501e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.539517796e-08 wvth0=1.549871091e-07 pvth0=-2.847194094e-14 k1=3.066737744e-01 lk1=9.013939151e-08 wk1=-3.067532285e-07 pk1=7.405762289e-14 k2=3.953484017e-02 lk2=-2.303623270e-08 wk2=6.211228500e-08 pk2=-1.743583257e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.997704092e-01 ldsub=4.205412629e-08 wdsub=-9.482212631e-07 pdsub=1.205429016e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.047939655e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.164255551e-09 wvoff=-1.608870732e-07 pvoff=2.958262129e-14 nfactor=3.512260001e+00 lnfactor=-2.877832618e-07 wnfactor=-4.353940989e-06 pnfactor=1.547337123e-12 eta0=0.49 etab=-2.667329801e-04 letab=-2.068124671e-11 wetab=2.943660666e-09 petab=-1.330184326e-15 u0=2.430190821e-02 lu0=-9.680288569e-10 wu0=1.994440090e-08 pu0=-5.570913243e-15 ua=-1.390389179e-09 lua=-1.582627219e-16 wua=1.472260752e-15 pua=-2.355837030e-22 ub=2.084225575e-18 lub=1.423312343e-25 wub=-6.607707533e-25 pub=-8.574311734e-32 uc=1.217486023e-11 luc=3.326293430e-17 wuc=4.837150578e-16 puc=-2.281862077e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.155206778e+04 lvsat=1.373292742e-02 wvsat=2.579412038e-01 pvsat=-5.972566178e-8 a0=1.5 ags=2.243633754e+00 lags=-4.490042142e-07 wags=-3.534518996e-12 pags=1.597181979e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.695053569e-02 lketa=-5.482500520e-09 wketa=6.688252317e-08 pketa=8.476717527e-15 dwg=0.0 dwb=0.0 pclm=1.173784523e+00 lpclm=-1.605465451e-07 wpclm=-3.756622035e-06 ppclm=8.056824773e-13 pdiblc1=3.031515126e+00 lpdiblc1=-7.806930142e-07 wpdiblc1=-9.237584483e-06 ppdiblc1=3.212936884e-12 pdiblc2=6.038826344e-03 lpdiblc2=-7.024633031e-10 wpdiblc2=-1.329185759e-08 ppdiblc2=2.655935385e-15 pdiblcb=5.403735547e-01 lpdiblcb=-2.554815673e-07 wpdiblcb=-2.827615197e-06 ppdiblcb=1.277745583e-12 drout=-1.797729302e+00 ldrout=5.648083892e-07 wdrout=1.324448636e-05 pdrout=-2.673810151e-12 pscbe1=-7.134173196e+08 lpscbe1=3.055302019e+02 wpscbe1=7.569087336e+03 ppscbe1=-1.528054920e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.945368856e-05 lalpha0=-8.370979114e-12 walpha0=-2.152234942e-10 palpha0=5.002373957e-17 alpha1=0.85 beta0=4.142412146e+01 lbeta0=-4.641204733e-06 wbeta0=-1.602475308e-04 pbeta0=3.332999353e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.202035728e-01 lkt1=-2.356337488e-08 wkt1=-3.115910144e-07 pkt1=1.268772615e-13 kt2=-4.498766624e-03 lkt2=-1.397989680e-08 wkt2=-1.991975655e-07 pkt2=8.798230898e-14 at=7.631297650e+04 lat=-1.080905910e-02 wat=-4.727104584e-03 pat=5.411118380e-9 ute=-1.217706545e+00 lute=-4.415653959e-08 wute=-4.622008321e-06 pute=1.735280338e-12 ua1=1.711277101e-09 lua1=-1.646676422e-16 wua1=-6.031228421e-15 pua1=2.016003981e-21 ub1=-2.027576640e-18 lub1=3.037017639e-25 wub1=3.356852845e-24 pub1=-1.022689421e-30 uc1=-1.232373589e-10 luc1=4.839997704e-17 wuc1=1.799740022e-16 puc1=-7.370939250e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.16 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.978392309e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.697884977e-08 wvth0=4.901940773e-07 pvth0=-9.614385887e-14 k1=5.037303652e-01 lk1=5.035740989e-08 wk1=1.580161711e-07 pk1=-1.977048828e-14 k2=-1.305220392e-02 lk2=-1.241990765e-08 wk2=-1.532207420e-07 pk2=2.603581425e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=9.847034013e-01 ldsub=-7.603273109e-08 wdsub=-8.908057895e-07 pdsub=1.089518084e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-7.267523460e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.364841706e-08 wvoff=-3.224256090e-07 pvoff=6.219418243e-14 nfactor=1.072634205e+00 lnfactor=2.047308337e-07 wnfactor=3.303890503e-06 pnfactor=1.366444095e-15 eta0=1.385914092e+00 leta0=-1.808680328e-07 weta0=-2.178746389e-07 peta0=4.398474998e-14 etab=6.725605415e-02 letab=-1.365224904e-08 wetab=-1.147963306e-07 petab=2.243928285e-14 u0=-2.439292397e-03 lu0=4.430511463e-09 wu0=2.656883467e-08 pu0=-6.908260557e-15 ua=-4.788360716e-09 lua=5.277231699e-16 wua=-1.728447067e-17 pua=6.512717610e-23 ub=4.370715641e-18 lub=-3.192676668e-25 wub=2.545188647e-24 pub=-7.329654070e-31 uc=3.237047706e-10 luc=-2.962903554e-17 wuc=-1.698021666e-15 puc=2.122649839e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.444451203e+04 lvsat=1.314899789e-02 wvsat=2.907268296e-01 pvsat=-6.634445671e-8 a0=1.5 ags=-2.298691977e+00 lags=4.680050466e-07 wags=1.262328213e-11 pags=-1.664771071e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.046308327e-01 lketa=1.019967552e-08 wketa=4.716553521e-07 pketa=-7.323922596e-14 dwg=0.0 dwb=0.0 pclm=1.055545655e+00 lpclm=-1.366763640e-07 wpclm=-2.849529799e-06 ppclm=6.225577896e-13 pdiblc1=-3.113588162e+00 lpdiblc1=4.598865826e-07 wpdiblc1=1.924023681e-05 ppdiblc1=-2.536194156e-12 pdiblc2=-7.072154243e-03 lpdiblc2=1.944394569e-09 wpdiblc2=-1.566805053e-08 ppdiblc2=3.135643591e-15 pdiblcb=-2.022045240e+00 lpdiblcb=2.618221015e-07 wpdiblcb=1.075289768e-05 ppdiblcb=-1.463901937e-12 drout=1.938809575e+00 ldrout=-1.895278158e-07 wdrout=-2.838671303e-06 pdrout=5.730738013e-13 pscbe1=8.156720299e+08 lpscbe1=-3.163885067e+00 wpscbe1=-5.559720697e+01 ppscbe1=1.122401974e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.260955972e-06 lalpha0=-8.624730672e-13 walpha0=3.734767448e-11 palpha0=-9.655805391e-19 alpha1=-2.241231372e+00 lalpha1=6.240608806e-07 walpha1=1.714339573e-05 palpha1=-3.460925874e-12 beta0=4.088528432e+01 lbeta0=-4.532423754e-06 wbeta0=-9.789918704e-05 pbeta0=2.074304754e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-5.480246079e-01 lkt1=4.261746351e-08 wkt1=1.365740805e-06 pkt1=-2.117441636e-13 kt2=-1.435019405e-01 lkt2=1.408220296e-08 wkt2=6.749977787e-07 pkt2=-8.850112129e-14 at=3.629549228e+04 lat=-2.730289368e-03 wat=-2.050713336e-01 pat=4.585681169e-8 ute=-7.492891382e-01 lute=-1.387211141e-07 wute=1.176707777e-05 pute=-1.573364751e-12 ua1=3.693450138e-09 lua1=-5.648307172e-16 wua1=1.095133633e-14 pua1=-1.412453173e-21 ub1=-3.873204422e-18 lub1=6.762989461e-25 wub1=-4.720408357e-25 pub1=-2.497085354e-31 uc1=-6.585054248e-11 luc1=3.681466915e-17 wuc1=5.433060218e-16 puc1=-1.470592240e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.17 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.734000131e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.676812847e-10 wvth0=8.849214844e-07 pvth0=-1.482009041e-13 k1=8.183162910e-01 lk1=8.869503414e-09 wk1=9.849192464e-08 pk1=-1.192037113e-14 k2=-6.259135231e-02 lk2=-5.886635220e-09 wk2=-4.238234297e-07 pk2=6.172316732e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.246663324e+00 ldsub=-1.105802677e-07 wdsub=-4.213465287e-06 pdsub=5.471474656e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=5.308807126e-02 lcdscd=-6.289149826e-09 wcdscd=-2.054852017e-07 pcdscd=2.709959388e-14 cit=0.0 voff='4.173915349e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.827891269e-08 wvoff=-2.508583719e-06 pvoff=3.505069001e-13 nfactor=1.872238091e+01 lnfactor=-2.122935412e-06 wnfactor=-8.002854834e-05 pnfactor=1.099133181e-11 eta0=6.035539042e-02 leta0=-6.052025680e-09 weta0=5.124328904e-07 peta0=-5.232893729e-14 etab=2.137548876e-02 letab=-7.601474191e-09 wetab=-9.842536475e-09 petab=8.597871528e-15 u0=5.133460555e-02 lu0=-2.661243972e-09 wu0=1.144358997e-07 pu0=-1.849625696e-14 ua=4.894456901e-09 lua=-7.492565002e-16 wua=4.218831777e-16 pua=7.209307470e-24 ub=-4.662166929e-18 lub=8.719979194e-25 wub=9.717682004e-24 pub=-1.678881003e-30 uc=1.576613818e-10 luc=-7.731067378e-18 wuc=2.921444656e-16 puc=-5.020011575e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.826274079e+05 lvsat=-2.437080598e-03 wvsat=-6.588027549e-01 pvsat=5.888045442e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.887311273e-01 lketa=1.136076065e-07 wketa=4.479320275e-06 pketa=-6.017740836e-13 dwg=0.0 dwb=0.0 pclm=-7.120591392e-01 lpclm=9.643712378e-08 wpclm=9.771193952e-06 ppclm=-1.041875879e-12 pdiblc1=-3.493929199e-02 lpdiblc1=5.387129101e-08 wpdiblc1=2.587828926e-06 ppdiblc1=-3.400579522e-13 pdiblc2=-4.196321082e-03 lpdiblc2=1.565126816e-09 wpdiblc2=7.402176466e-08 ppdiblc2=-8.692738926e-15 pdiblcb=-4.656752491e-01 lpdiblcb=5.656647069e-08 wpdiblcb=6.026978841e-07 ppdiblcb=-1.252834380e-13 drout=-1.170919074e-01 ldrout=8.160652760e-08 wdrout=1.012642254e-05 pdrout=-1.136775740e-12 pscbe1=8.099807356e+08 lpscbe1=-2.413311486e+00 wpscbe1=2.885653283e+01 ppscbe1=8.617608125e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.891174542e-05 lalpha0=1.929803965e-12 walpha0=1.319956040e-10 palpha0=-1.344784413e-17 alpha1=8.062873201e+00 lalpha1=-7.348547346e-07 walpha1=-4.000125671e-05 palpha1=4.075368035e-12 beta0=-1.841674107e+01 lbeta0=3.288386657e-06 wbeta0=2.610668285e-04 pbeta0=-2.659774955e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.694683401e-01 lkt1=3.225738436e-08 wkt1=4.334108265e-07 pkt1=-8.878755368e-14 kt2=-5.934223412e-02 lkt2=2.983136714e-09 wkt2=2.339152909e-09 pkt2=2.097709304e-16 at=1.788698181e+05 lat=-2.153313403e-02 wat=-9.235371282e-01 pat=1.406087991e-7 ute=-7.917937163e+00 lute=8.066873562e-07 wute=-7.170255859e-07 pute=7.305128372e-14 ua1=-1.079852373e-08 lua1=1.346385289e-15 wua1=1.130248717e-14 pua1=-1.458763297e-21 ub1=6.735780990e-18 lub1=-7.228246591e-25 wub1=-6.115646489e-24 pub1=4.945758218e-31 uc1=2.397279496e-10 luc1=-3.485327963e-18 wuc1=-1.403030367e-15 puc1=1.096255653e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.18 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.235866060e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.285945491e-07 wvth0=-6.759846982e-09 pvth0=6.756594211e-13 k1=5.438745012e-01 lk1=-3.007403405e-07 wk1=-1.696621638e-08 pk1=1.695805240e-12 k2=-2.823294061e-02 lk2=1.419266340e-07 wk2=5.607470331e-09 pk2=-5.604772073e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.061890569e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.200140101e-08 wvoff=3.121632721e-09 pvoff=-3.120130623e-13 nfactor=2.513979061e+00 lnfactor=6.787826135e-06 wnfactor=-3.144637240e-08 pnfactor=3.143124072e-12 eta0=0.08 etab=-0.07 u0=3.239173954e-02 lu0=-1.300328259e-09 wu0=1.037355928e-09 pu0=-1.036856762e-13 ua=-7.622581428e-10 lua=2.645199369e-16 wua=-3.360801101e-17 pua=3.359183918e-21 ub=1.749717917e-18 lub=-1.388453243e-24 wub=6.463352613e-26 pub=-6.460242513e-30 uc=5.890830949e-11 luc=-9.661658154e-16 wuc=-4.527716083e-17 puc=4.525537392e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.312864498e+00 la0=-1.592083312e-06 wa0=-1.222009775e-07 pa0=1.221421756e-11 ags=4.457152188e-01 lags=-9.241769639e-07 wags=-3.263253706e-08 pags=3.261683460e-12 a1=0.0 a2=0.42385546 b0=7.886836216e-25 lb0=-7.883041149e-29 wb0=-3.944460748e-30 pb0=3.942562713e-34 b1=2.632910460e-24 lb1=-5.253151618e-29 keta=-9.246939892e-03 lketa=4.521222310e-08 wketa=-9.902814569e-10 pketa=9.898049434e-14 dwg=0.0 dwb=0.0 pclm=1.619338699e-02 lpclm=1.011774211e-06 wpclm=-1.244565060e-08 ppclm=1.243966188e-12 pdiblc1=0.39 pdiblc2=2.769830753e-03 lpdiblc2=3.034818446e-08 wpdiblc2=1.368575327e-09 ppdiblc2=-1.367916782e-13 pdiblcb=-9.556476466e-01 lpdiblcb=9.301998282e-05 wpdiblcb=4.654468549e-06 ppdiblcb=-4.652228865e-10 drout=0.56 pscbe1=8.067205144e+08 lpscbe1=-5.202131024e+03 wpscbe1=-1.852818016e+02 ppscbe1=1.851926458e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.071777822e-01 lkt1=-5.849401785e-07 wkt1=-1.508677152e-08 pkt1=1.507951192e-12 kt2=-4.359975286e-02 lkt2=-1.712759580e-07 wkt2=-8.325503837e-09 pkt2=8.321497688e-13 at=140000.0 ute=-1.760911156e+00 lute=-5.246358714e-06 wute=-1.748268561e-07 pute=1.747427312e-11 ua1=4.320442450e-10 lua1=-5.599728672e-15 wua1=-1.343583697e-16 pua1=1.342937178e-20 ub1=-6.477720772e-19 lub1=8.148154486e-25 wub1=-1.360617149e-25 pub1=1.359962433e-29 uc1=1.483515271e-11 luc1=9.940817173e-17 wuc1=3.480804577e-18 puc1=-3.479129648e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.19 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.121293129e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.710460024e-8 k1=5.288012186e-01 wk1=6.802853878e-8 k2=-2.111949431e-02 wk2=-2.248397665e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.015778926e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.251664531e-8 nfactor=2.854188895e+00 wnfactor=1.260888531e-7 eta0=0.08 etab=-0.07 u0=3.232656633e-02 wu0=-4.159431094e-9 ua=-7.490002481e-10 wua=1.347562609e-16 ub=1.680127824e-18 wub=-2.591576248e-25 uc=1.048351107e-11 wuc=1.815454326e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.233068347e+00 wa0=4.899827841e-7 ags=3.993949263e-01 wags=1.308449546e-7 a1=0.0 a2=0.42385546 b0=-3.162342925e-24 wb0=1.581589524e-29 b1=0.0 keta=-6.980876703e-03 wketa=3.970679083e-9 dwg=0.0 dwb=0.0 pclm=6.690410501e-02 wpclm=4.990266572e-8 pdiblc1=0.39 pdiblc2=4.290899591e-03 wpdiblc2=-5.487503969e-9 pdiblcb=3.706568554e+00 wpdiblcb=-1.866277590e-5 drout=0.56 pscbe1=5.459866506e+08 wpscbe1=7.429146217e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.364953277e-01 wkt1=6.049262832e-8 kt2=-5.218420452e-02 wkt2=3.338233157e-8 at=140000.0 ute=-2.023861737e+00 wute=7.009939808e-7 ua1=1.513825534e-10 wua1=5.387296354e-16 ub1=-6.069330481e-19 wub1=5.455594482e-25 uc1=1.981754869e-11 wuc1=-1.395679766e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.20 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.967908026e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.219700082e-07 wvth0=6.048249080e-08 pvth0=-2.654170138e-13 k1=5.141396921e-01 lk1=1.165867145e-07 wk1=1.026764709e-07 pk1=-2.755162332e-13 k2=-9.542306900e-03 lk2=-9.206041659e-08 wk2=-4.545107818e-08 pk2=1.826316583e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016409368e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.013198553e-10 wvoff=-1.838554534e-08 pvoff=4.666879465e-14 nfactor=3.804650792e+00 lnfactor=-7.557959896e-06 wnfactor=-3.350731493e-06 pnfactor=2.764726165e-11 eta0=0.08 etab=-0.07 u0=3.031615667e-02 lu0=1.598653832e-08 wu0=3.007168460e-09 pu0=-5.698794683e-14 ua=-6.441389313e-10 lua=-8.338447134e-16 wua=-3.415772470e-16 pua=3.787747371e-21 ub=1.335116414e-18 lub=2.743489677e-24 wub=1.057227702e-24 pub=-1.046773947e-29 uc=-1.032858754e-10 luc=9.046806225e-16 wuc=5.536228242e-16 puc=-2.958715141e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=9.752769239e-01 la0=2.049926716e-06 wa0=1.722259742e-06 pa0=-9.798919730e-12 ags=2.390936052e-01 lags=1.274697030e-06 wags=5.810890742e-07 pags=-3.580287659e-12 a1=0.0 a2=0.42385546 b0=-6.286643656e-24 lb0=2.484406762e-29 wb0=3.144152922e-29 pb0=-1.242531819e-34 b1=0.0 keta=-9.951967801e-03 lketa=2.362576286e-08 wketa=-1.853873304e-09 pketa=4.631614746e-14 dwg=0.0 dwb=0.0 pclm=-3.534741081e-01 lpclm=3.342797525e-06 wpclm=1.097343179e-07 ppclm=-4.757741779e-13 pdiblc1=0.39 pdiblc2=5.717396704e-03 lpdiblc2=-1.134333529e-08 wpdiblc2=-1.281910512e-08 ppdiblc2=5.830001986e-14 pdiblcb=7.393247270e+00 lpdiblcb=-2.931603044e-05 wpdiblcb=-3.710104327e-05 ppdiblcb=1.466189080e-10 drout=0.56 pscbe1=2.976693751e+08 lpscbe1=1.974589425e+03 wpscbe1=1.468967605e+03 ppscbe1=-5.773486924e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.577231195e-01 lkt1=1.688008748e-07 wkt1=1.307868485e-07 pkt1=-5.589712736e-13 kt2=-6.264076055e-02 lkt2=8.314928920e-08 wkt2=6.802786124e-08 pkt2=-2.754971291e-13 at=140000.0 ute=-2.366573280e+00 lute=2.725201402e-06 wute=1.648631252e-06 pute=-7.535498815e-12 ua1=-4.886511121e-10 lua1=5.089471544e-15 wua1=2.590875593e-15 pua1=-1.631842045e-20 ub1=-1.849308792e-19 lub1=-3.355711029e-24 wub1=-9.416822838e-25 pub1=1.182636927e-29 uc1=2.793341020e-11 luc1=-6.453636491e-17 wuc1=-7.384980154e-17 puc1=4.762620395e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.21 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.284356918e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.086828136e-09 wvth0=-3.282894099e-08 pvth0=1.033386606e-13 k1=5.393792916e-01 lk1=1.684282089e-08 wk1=3.201483368e-09 pk1=1.175970800e-13 k2=-3.056306260e-02 lk2=-8.988891525e-09 wk2=1.695146791e-08 pk2=-6.397577797e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.292148904e+00 ldsub=-2.893365343e-06 wdsub=-2.197414613e-06 pdsub=8.683921058e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064940750e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.968034423e-08 wvoff=2.286693560e-10 pvoff=-2.689236673e-14 nfactor=1.080033482e+00 lnfactor=3.209403481e-06 wnfactor=6.874124785e-06 pnfactor=-1.276015360e-11 eta0=2.740194596e-01 leta0=-7.667418159e-07 weta0=-5.823148724e-07 peta0=2.301239080e-12 etab=-2.396144958e-01 letab=6.702963034e-07 wetab=5.090677178e-07 petab=-2.011775042e-12 u0=3.785839604e-02 lu0=-1.381949414e-08 wu0=-2.082848193e-08 pu0=3.720770709e-14 ua=-8.781557840e-10 lua=9.096204051e-17 wua=1.114086925e-15 pua=-1.964864214e-21 ub=2.366368951e-18 lub=-1.331897630e-24 wub=-3.203067539e-24 pub=6.368440347e-30 uc=1.668307468e-10 luc=-1.627881244e-16 wuc=-3.288410595e-16 puc=5.286771140e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.326372002e+00 la0=-3.289440253e-06 wa0=-4.023470549e-06 pa0=1.290752264e-11 ags=6.306909225e-01 lags=-2.728489683e-07 wags=-1.245143297e-06 pags=3.636765352e-12 a1=0.0 a2=0.42385546 b0=3.086258536e-24 lb0=-1.219652647e-29 wb0=-1.543537271e-29 pb0=6.099875615e-35 b1=0.0 keta=-1.066419448e-02 lketa=2.644039792e-08 wketa=2.679651307e-08 pketa=-6.690677008e-14 dwg=0.0 dwb=0.0 pclm=6.021686271e-01 lpclm=-4.337888424e-07 wpclm=-3.846574773e-07 ppclm=1.478003364e-12 pdiblc1=0.39 pdiblc2=3.390211118e-04 lpdiblc2=9.911365026e-09 wpdiblc2=5.483873308e-09 ppdiblc2=-1.403117281e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.825068970e+08 lpscbe1=5.856923401e+01 wpscbe1=7.692721352e+01 ppscbe1=-2.723089492e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.954274373e-01 lkt1=-7.738424810e-08 wkt1=-5.900063168e-08 pkt1=1.910462633e-13 kt2=-4.018570198e-02 lkt2=-5.590430100e-09 wkt2=-7.534194070e-09 pkt2=2.311512159e-14 at=1.616895874e+05 lat=-8.571466818e-02 wat=7.837445453e-03 pat=-3.097265177e-8 ute=-1.520398050e+00 lute=-6.187824119e-07 wute=-1.247750985e-06 pute=3.910659116e-12 ua1=1.253832652e-09 lua1=-1.796616937e-15 wua1=-3.665691139e-15 pua1=8.406786743e-21 ub1=-1.506908123e-18 lub1=1.868585723e-24 wub1=3.637091864e-24 pub1=-6.268401287e-30 uc1=3.213453451e-12 luc1=3.315396248e-17 wuc1=1.995144897e-17 puc1=1.055706599e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.22 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.127695596e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.749159764e-08 wvth0=-4.451959181e-08 pvth0=1.261574198e-13 k1=4.334189857e-01 lk1=2.236647287e-07 wk1=5.862048552e-07 pk1=-1.020356124e-12 k2=4.127113612e-03 lk2=-7.669998736e-08 wk2=-1.949083613e-07 pk2=3.495493974e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.477883764e+00 ldsub=2.513408792e-06 wdsub=6.973415792e-06 pdsub=-9.216448563e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.549663687e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.130415623e-08 wvoff=4.753663013e-08 pvoff=-1.192318765e-13 nfactor=2.556902913e+00 lnfactor=3.267301006e-07 wnfactor=2.400182664e-06 pnfactor=-4.027550980e-12 eta0=-2.294484072e-01 leta0=2.159675473e-07 weta0=1.150074892e-06 peta0=-1.080179585e-12 etab=8.308667538e-02 letab=4.042201862e-08 wetab=-4.183944493e-07 petab=-2.014792596e-13 u0=3.457069975e-02 lu0=-7.402302221e-09 wu0=-4.461785572e-10 pu0=-2.576123608e-15 ua=-3.601346315e-10 lua=-9.201536047e-16 wua=6.513555324e-16 pua=-1.061667600e-21 ub=1.218455784e-18 lub=9.086922703e-25 wub=-3.288606877e-25 pub=7.583306035e-31 uc=1.494617889e-10 luc=-1.288859856e-16 wuc=-2.869198883e-16 puc=4.468519766e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.448626720e+04 lvsat=3.028096029e-02 wvsat=5.917492718e-02 pvsat=-1.155024160e-7 a0=-7.488554919e-01 la0=2.713037863e-06 wa0=8.361131609e-06 pa0=-1.126574701e-11 ags=-5.068486146e-01 lags=1.947492841e-06 wags=2.291367490e-06 pags=-3.266082861e-12 a1=0.0 a2=0.42385546 b0=-6.172517071e-24 lb0=5.875501722e-30 wb0=3.087074542e-29 pb0=-2.938527603e-35 b1=0.0 keta=9.155753608e-02 lketa=-1.730842557e-07 wketa=-1.259120035e-07 pketa=2.311620820e-13 dwg=0.0 dwb=0.0 pclm=1.215939487e+00 lpclm=-1.631796522e-06 wpclm=-3.236943703e-06 ppclm=7.045326655e-12 pdiblc1=2.289559520e-01 lpdiblc1=3.143388175e-07 wpdiblc1=-1.753706799e-07 ppdiblc1=3.423026980e-13 pdiblc2=3.238907380e-03 lpdiblc2=4.251132118e-09 wpdiblc2=9.314340086e-09 ppdiblc2=-2.150778814e-14 pdiblcb=-4.884024301e-02 lpdiblcb=4.653331737e-08 wpdiblcb=6.773034642e-10 ppdiblcb=-1.322015763e-15 drout=8.455643000e-01 ldrout=-5.573875314e-7 pscbe1=5.791628579e+08 lpscbe1=4.554726004e+02 wpscbe1=1.700416500e+03 ppscbe1=-3.441166842e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.997924372e-06 lalpha0=1.762143405e-11 walpha0=2.701342927e-11 palpha0=-5.272699934e-17 alpha1=1.084756326e+00 lalpha1=-4.582164117e-07 walpha1=-1.335954531e-06 palpha1=2.607624266e-12 beta0=7.558002181e+00 lbeta0=1.230074981e-05 wbeta0=1.700305767e-05 pbeta0=-3.318794521e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.669878830e-01 lkt1=6.229322613e-08 wkt1=-5.723510189e-08 pkt1=1.876001592e-13 kt2=-7.230996607e-02 lkt2=5.711231061e-08 wkt2=7.560597679e-08 pkt2=-1.391645982e-13 at=1.757976144e+05 lat=-1.132518581e-01 wat=-4.084217390e-02 pat=6.404417232e-8 ute=-3.251468453e+00 lute=2.760061018e-06 wute=3.822478576e-06 pute=-5.985825628e-12 ua1=-2.478219363e-09 lua1=5.487904484e-15 wua1=5.973869460e-15 pua1=-1.040848844e-20 ub1=5.166393454e-19 lub1=-2.081138133e-24 wub1=2.004958755e-25 pub1=4.394251280e-31 uc1=-1.027501739e-10 luc1=2.399823535e-16 wuc1=6.146364423e-16 puc1=-1.055183680e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.23 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.042618932e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.558988367e-08 wvth0=2.069055047e-07 pvth0=-1.131693525e-13 k1=9.759198267e-01 lk1=-2.927315143e-07 wk1=-1.600327074e-06 pk1=1.060962075e-12 k2=-1.843737641e-01 lk2=1.027304166e-07 wk2=5.527076651e-07 pk2=-3.620920934e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.854795310e+00 ldsub=-6.589050976e-07 wdsub=-4.976018670e-06 pdsub=2.157991062e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-7.868648734e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.778660818e-08 wvoff=-1.499990683e-07 pvoff=6.879860168e-14 nfactor=3.160238432e+00 lnfactor=-2.475735171e-07 wnfactor=-3.834408655e-06 pnfactor=1.907038039e-12 eta0=-4.477234439e-01 leta0=4.237394075e-07 weta0=2.910970639e-08 peta0=-1.315412323e-14 etab=2.388798930e-01 letab=-1.078745852e-07 wetab=-1.197362287e-06 petab=5.400054246e-13 u0=2.809610460e-02 lu0=-1.239258113e-09 wu0=1.551945934e-09 pu0=-4.478100347e-15 ua=-1.182123076e-09 lua=-1.377184219e-16 wua=-5.958541054e-16 pua=1.255275572e-22 ub=2.141486556e-18 lub=3.007681594e-26 wub=7.952333845e-25 pub=-3.116731860e-31 uc=-5.469178900e-11 luc=6.544392635e-17 wuc=3.863433334e-16 puc=-1.940144922e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.082429701e+04 lvsat=1.472910014e-02 wvsat=-1.349410598e-01 pvsat=6.927290381e-8 a0=2.644790098e+00 la0=-5.173088941e-07 wa0=-6.613889380e-06 pa0=2.988690947e-12 ags=1.711394680e+00 lags=-1.640108049e-07 wags=-1.724982902e-06 pags=5.570047664e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.704751193e-01 lketa=7.633965031e-08 wketa=3.149244014e-07 pketa=-1.884617159e-13 dwg=0.0 dwb=0.0 pclm=-1.364184711e+00 lpclm=8.241746800e-07 wpclm=8.090192979e-06 ppclm=-3.736759537e-12 pdiblc1=-2.427067727e-01 lpdiblc1=7.633056035e-07 wpdiblc1=2.918015320e-06 ppdiblc1=-2.602232661e-12 pdiblc2=9.367445421e-03 lpdiblc2=-1.582506801e-09 wpdiblc2=-1.233987224e-08 ppdiblc2=-8.955548576e-16 pdiblcb=2.268048603e-02 lpdiblcb=-2.154590571e-08 wpdiblcb=-1.354606928e-09 ppdiblcb=6.121211334e-16 drout=-2.218191936e-01 ldrout=4.586345358e-07 wdrout=-5.611412266e-07 pdrout=5.341396720e-13 pscbe1=1.290523841e+09 lpscbe1=-2.216584040e+02 wpscbe1=-3.645145366e+03 ppscbe1=1.647171933e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.243938038e-05 lalpha0=-1.230313904e-11 walpha0=-7.580027212e-11 palpha0=4.513940955e-17 alpha1=3.804873487e-01 lalpha1=2.121638464e-07 walpha1=2.671909063e-06 palpha1=-1.207384939e-12 beta0=3.210324317e+01 lbeta0=-1.106339873e-05 wbeta0=-6.220980807e-05 pbeta0=4.221327664e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.232778930e-01 lkt1=2.068651717e-08 wkt1=2.708073996e-07 pkt1=-1.246572651e-13 kt2=8.604100608e-03 lkt2=-1.990825210e-08 wkt2=-1.304050438e-07 pkt2=5.693337808e-14 at=4.968215630e+04 lat=6.795050241e-03 wat=9.950071098e-02 pat=-6.954555328e-8 ute=9.568367684e-01 lute=-1.245744765e-06 wute=-6.178040085e-06 pute=3.533478075e-12 ua1=5.336087769e-09 lua1=-1.950386004e-15 wua1=-9.503107640e-15 pua1=4.323752001e-21 ub1=-1.394890363e-18 lub1=-2.615893226e-25 wub1=-2.522531016e-24 pub1=3.031422689e-30 uc1=3.837568618e-10 luc1=-2.231144503e-16 wuc1=-1.379726595e-15 puc1=8.432126028e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.24 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.336652932e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.288505416e-08 wvth0=-6.342383903e-08 pvth0=8.987341660e-15 k1=-8.210769466e-03 lk1=1.519784036e-07 wk1=1.268085768e-06 pk1=-2.352191886e-13 k2=1.376072839e-01 lk2=-4.276670135e-08 wk2=-4.283795853e-07 pk2=8.124259436e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.257618329e-01 ldsub=3.203607887e-08 wdsub=-5.780805422e-07 pdsub=1.706463826e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.400773430e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.524695099e-11 wvoff=1.557645867e-08 pvoff=-6.021833043e-15 nfactor=2.697206512e+00 lnfactor=-3.833819003e-08 wnfactor=-2.775960411e-07 pnfactor=2.997819984e-13 eta0=0.49 etab=1.742734697e-03 letab=-7.168089498e-10 wetab=-7.106334237e-09 petab=2.151374471e-15 u0=3.071902501e-02 lu0=-2.424506009e-09 wu0=-1.214966650e-08 pu0=1.713397980e-15 ua=-9.509803612e-10 lua=-2.421674231e-16 wua=-7.253642364e-16 pua=1.840507247e-22 ub=1.854110405e-18 lub=1.599366386e-25 wub=4.901093082e-25 pub=-1.737934133e-31 uc=1.568570550e-10 luc=-3.015097682e-17 wuc=-2.398871859e-16 puc=8.896718109e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.219547645e+05 lvsat=-3.856976660e-03 wvsat=-4.415213242e-02 pvsat=2.824711249e-8 a0=1.5 ags=2.421571483e+00 lags=-4.849262085e-07 wags=-8.899274135e-07 pags=1.796590574e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.414948712e-02 lketa=-7.088701473e-09 wketa=-1.386719251e-07 pketa=1.650984569e-14 dwg=0.0 dwb=0.0 pclm=3.613279008e-01 lpclm=4.444831533e-08 wpclm=3.067351451e-07 ppclm=-2.195628281e-13 pdiblc1=1.794079288e+00 lpdiblc1=-1.570793184e-07 wpdiblc1=-3.048769405e-06 ppdiblc1=9.404398746e-14 pdiblc2=8.616990966e-03 lpdiblc2=-1.243390692e-09 wpdiblc2=-2.618608904e-08 ppdiblc2=5.361287436e-15 pdiblcb=-2.673639547e-01 lpdiblcb=1.095196662e-07 wpdiblcb=1.212140179e-06 ppdiblcb=-5.477431160e-13 drout=6.260706271e-01 ldrout=7.548923573e-08 wdrout=1.122282453e-06 pdrout=-2.265675040e-13 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.374087929e-05 lalpha0=4.046032884e-12 walpha0=5.081966822e-11 palpha0=-1.207773571e-17 alpha1=0.85 beta0=-2.231082189e+00 lbeta0=4.451630547e-06 wbeta0=5.808619960e-05 pbeta0=-1.214620360e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.476669907e-01 lkt1=-1.348061298e-08 wkt1=-1.742376182e-07 pkt1=7.645012254e-14 kt2=-3.143232691e-02 lkt2=-1.816551193e-09 wkt2=-6.449415788e-08 pkt2=2.714950102e-14 at=8.958442304e+04 lat=-1.123602595e-02 wat=-7.110188210e-02 pat=7.546517087e-9 ute=-2.297161941e+00 lute=2.246754258e-07 wute=7.766956977e-07 pute=3.907651151e-13 ua1=1.332413964e-09 lua1=-1.412018811e-16 wua1=-4.136411880e-15 pua1=1.898644154e-21 ub1=-3.571200901e-18 lub1=7.218440597e-25 wub1=1.107701482e-23 pub1=-3.113953684e-30 uc1=-2.978064402e-10 luc1=8.487105622e-17 wuc1=1.053050189e-15 puc1=-2.561130032e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.25 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='7.892227260e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.428914423e-08 wvth0=-4.669764070e-07 pvth0=9.045693763e-14 k1=5.321744500e-01 lk1=4.288489509e-08 wk1=1.575814439e-08 pk1=1.760196434e-14 k2=-5.423093901e-02 lk2=-4.038209072e-09 wk2=5.272737177e-08 pk2=-1.588375924e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.317057938e-01 ldsub=-7.010439391e-08 wdsub=-1.256154893e-07 pdsub=7.930228524e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-4.065689119e-03 lcdscd=1.910942785e-09 wcdscd=4.734095924e-08 pcdscd=-9.557240192e-15 cit=0.0 voff='-2.298582160e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.807980549e-08 wvoff=4.636970940e-07 pvoff=-9.648887502e-14 nfactor=-1.576788206e+00 lnfactor=8.245001375e-07 wnfactor=1.655450509e-05 pnfactor=-3.098299410e-12 eta0=1.238041915e+00 leta0=-1.510154499e-07 weta0=5.216817319e-07 peta0=-1.053176297e-13 etab=-3.115441362e-02 letab=5.924500250e-09 wetab=3.773861069e-07 petab=-7.547034404e-14 u0=8.285319580e-03 lu0=2.104432876e-09 wu0=-2.706840315e-08 pu0=4.725207455e-15 ua=-6.229252515e-09 lua=8.234154375e-16 wua=7.189079382e-15 pua=-1.413725067e-21 ub=7.464087282e-18 lub=-9.726111034e-25 wub=-1.292575900e-23 pub=2.534615496e-30 uc=-1.926866093e-10 luc=4.041524768e-17 wuc=8.846179028e-16 puc=-1.380490307e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.962905475e+04 lvsat=6.501599590e-04 wvsat=1.147576020e-01 pvsat=-3.833743601e-9 a0=1.5 ags=-2.298688371e+00 lags=4.680045711e-07 wags=-5.411340083e-12 pags=7.136529417e-19 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.496907703e-03 lketa=-4.938148087e-09 wketa=-6.912629484e-08 pketa=2.469904302e-15 dwg=0.0 dwb=0.0 pclm=5.459899473e-01 lpclm=7.168556715e-09 wpclm=-3.010776299e-07 ppclm=-9.685697721e-14 pdiblc1=2.170773015e+00 lpdiblc1=-2.331266247e-07 wpdiblc1=-7.188555006e-06 ppdiblc1=9.297880443e-13 pdiblc2=-1.292503406e-02 lpdiblc2=3.105534861e-09 wpdiblc2=1.360408604e-08 ppdiblc2=-2.671592900e-15 pdiblcb=1.001738217e+00 lpdiblcb=-1.466879493e-07 wpdiblcb=-4.370017047e-06 ppdiblcb=5.791883668e-13 drout=5.240808131e-01 ldrout=9.607904136e-08 wdrout=4.236842777e-06 pdrout=-8.553380567e-13 pscbe1=7.871335424e+08 lpscbe1=2.597493333e+00 wpscbe1=8.713295853e+01 ppscbe1=-1.759048880e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.013037805e-05 lalpha0=-7.731204195e-13 walpha0=-2.009839292e-12 palpha0=-1.412461902e-18 alpha1=1.691576134e+00 lalpha1=-1.698982314e-07 walpha1=-2.525840964e-06 palpha1=5.099192997e-13 beta0=1.079891952e+01 lbeta0=1.821120772e-06 wbeta0=5.257241116e-05 pbeta0=-1.103307447e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.310243157e-01 lkt1=3.347647158e-09 wkt1=2.804524700e-07 pkt1=-1.534316714e-14 kt2=-2.894316139e-02 lkt2=-2.319066418e-09 wkt2=1.020524362e-07 pkt2=-6.473091949e-15 at=1.040979730e+05 lat=-1.416603594e-02 wat=-5.441733724e-01 pat=1.030506626e-7 ute=1.494709572e+00 lute=-5.408313870e-07 wute=5.441176509e-07 pute=4.377182038e-13 ua1=4.307800179e-09 lua1=-7.418758255e-16 wua1=7.878773956e-15 pua1=-5.269935777e-22 ub1=-1.670196568e-18 lub1=3.380674040e-25 wub1=-1.148999248e-23 pub1=1.441896317e-30 uc1=3.034084642e-10 luc1=-3.650280989e-17 wuc1=-1.303477172e-15 puc1=2.196250970e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.26 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.453990170e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.213342967e-08 wvth0=5.248312819e-07 pvth0=-4.034365218e-14 k1=7.343677863e-01 lk1=1.621943571e-08 wk1=5.183454282e-07 pk1=-4.867974923e-14 k2=-1.278931595e-01 lk2=5.676438230e-09 wk2=-9.722806478e-08 pk2=3.892513683e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.224763809e-01 ldsub=-2.946709694e-09 wdsub=4.086912039e-07 pdsub=8.837384240e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.693329888e-02 lcdscd=-2.177234751e-09 wcdscd=-7.467678971e-08 pcdscd=6.534582557e-15 cit=0.0 voff='6.264320214e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.049557404e-08 wvoff=-7.343730776e-07 pvoff=6.151381728e-14 nfactor=8.278561148e+00 lnfactor=-4.752331906e-07 wnfactor=-2.779564278e-05 pnfactor=2.750642441e-12 eta0=4.061031411e-01 leta0=-4.129853242e-08 weta0=-1.216762942e-06 peta0=1.239501923e-13 etab=1.253069003e-01 letab=-1.470977429e-08 wetab=-5.296369914e-07 petab=4.414876919e-14 u0=1.243356313e-01 lu0=-1.320039828e-08 wu0=-2.506657363e-07 pu0=3.421344734e-14 ua=1.432770838e-08 lua=-1.887657122e-15 wua=-4.675684499e-14 pua=5.700717384e-21 ub=-1.233392251e-17 lub=1.638370225e-24 wub=4.808660195e-23 pub=-5.511755677e-30 uc=4.506819141e-10 luc=-4.443283656e-17 wuc=-1.173345569e-15 puc=1.333572499e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.834607187e+04 lvsat=1.620883763e-02 wvsat=3.463303307e-01 pvsat=-3.437378664e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.458313643e-01 lketa=-6.327365856e-08 wketa=-2.195256475e-06 pketa=2.828660786e-13 dwg=0.0 dwb=0.0 pclm=2.233844459e+00 lpclm=-2.154273841e-07 wpclm=-4.962218522e-06 ppclm=5.178589448e-13 pdiblc1=6.708489545e-01 lpdiblc1=-3.531513965e-08 wpdiblc1=-9.420453585e-07 ppdiblc1=1.059921056e-13 pdiblc2=1.390258127e-02 lpdiblc2=-4.325178750e-10 wpdiblc2=-1.649667383e-08 ppdiblc2=1.298125414e-15 pdiblcb=-7.081350585e-01 lpdiblcb=7.881184814e-08 wpdiblcb=1.815317463e-06 ppdiblcb=-2.365397337e-13 drout=4.015081417e+00 ldrout=-3.643176092e-07 wdrout=-1.053990681e-05 pdrout=1.093434456e-12 pscbe1=8.522625542e+08 lpscbe1=-5.991785873e+00 wpscbe1=-1.826084565e+02 ppscbe1=1.798327876e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.866091795e-05 lalpha0=-1.898136551e-12 walpha0=-5.591738391e-11 palpha0=5.696918990e-18 alpha1=-1.113677645e+00 lalpha1=2.000614421e-07 walpha1=5.893628917e-06 palpha1=-6.004488077e-13 beta0=6.110741390e+01 lbeta0=-4.813613775e-06 wbeta0=-1.366590773e-04 pbeta0=1.392296345e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-5.806687605e-01 lkt1=3.627100618e-08 wkt1=9.895599357e-07 pkt1=-1.088609688e-13 kt2=-1.038877366e-01 lkt2=7.564699104e-09 wkt2=2.251255544e-07 pkt2=-2.270409784e-14 at=-2.045509893e+05 lat=2.653889786e-02 wat=9.940737912e-01 pat=-9.981491156e-8 ute=-1.817915277e+01 lute=2.053777253e-06 wute=5.060261778e-05 pute=-6.164046851e-12 ua1=-2.131641681e-08 lua1=2.637471535e-15 wua1=6.390585718e-14 pua1=-7.915901341e-21 ub1=1.272398400e-17 lub1=-1.560251524e-24 wub1=-3.606457795e-23 pub1=4.682817224e-30 uc1=-3.229135141e-10 luc1=4.609715893e-17 wuc1=1.410920764e-15 puc1=-1.383524172e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.27 nmos lmin=2.0e-05 lmax=0.0001 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.307128993e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.905943188e-07 wvth0=-2.814814772e-08 pvth0=5.616084937e-13 k1=5.343766968e-01 lk1=3.409918755e-07 wk1=1.153975295e-08 pk1=-2.302397777e-13 k2=-2.935986967e-02 lk2=1.494431142e-08 wk2=8.989747324e-09 pk2=-1.793623688e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.081196041e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.731257626e-08 wvoff=8.915826504e-09 pvoff=-1.778875094e-13 nfactor=1.759593052e+00 lnfactor=2.267744657e-05 wnfactor=2.232708952e-06 pnfactor=-4.454674332e-11 eta0=0.08 etab=-0.07 u0=3.494734414e-02 lu0=-7.994008717e-08 wu0=-6.632836385e-09 pu0=1.323375622e-13 ua=-8.673616060e-10 lua=3.257350596e-15 wua=2.818413253e-16 pua=-5.623264582e-21 ub=2.040092932e-18 lub=-8.904782501e-24 wub=-8.068753943e-25 pub=1.609868185e-29 uc=4.997117375e-11 luc=4.190059862e-16 wuc=-1.845393873e-17 puc=3.681907896e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.186875978e+00 la0=4.178882018e-06 wa0=2.559311397e-07 pa0=-5.106307644e-12 ags=4.621273943e-01 lags=-3.818130466e-07 wags=-8.189076025e-08 pags=1.633874704e-12 a1=0.0 a2=0.42385546 b0=-5.255574854e-25 lb0=5.253045924e-29 b1=7.902212087e-24 lb1=-1.576639952e-28 wb1=-1.581487090e-29 pb1=3.155364222e-34 keta=-1.609718144e-02 lketa=2.082833011e-07 wketa=1.956949922e-08 pketa=-3.904483196e-13 dwg=0.0 dwb=0.0 pclm=-1.143910264e-01 lpclm=3.948916717e-06 wpclm=3.794802220e-07 ppclm=-7.571344232e-12 pdiblc1=0.39 pdiblc2=2.925192138e-03 lpdiblc2=-9.230834263e-09 wpdiblc2=9.022857848e-10 ppdiblc2=-1.800229861e-14 pdiblcb=5.951584812e-01 lpdiblcb=-6.198600671e-05 wpdiblcb=-1.110223025e-22 ppdiblcb=-7.105427358e-27 drout=0.56 pscbe1=8.953737561e+08 lpscbe1=-2.032258218e+03 wpscbe1=-4.513587262e+02 ppscbe1=9.005455593e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.837743889e-01 lkt1=-6.497451980e-07 wkt1=-8.532789077e-08 pkt1=1.702451923e-12 kt2=-4.588319540e-02 lkt2=9.619866054e-08 wkt2=-1.472157522e-09 pkt2=2.937231168e-14 at=140000.0 ute=-1.643379560e+00 lute=-2.931339137e-06 wute=-5.275770203e-07 pute=1.052615393e-11 ua1=6.796303143e-10 lua1=-6.958224771e-15 wua1=-8.774438864e-16 pua1=1.750665601e-20 ub1=-1.047594621e-18 lub1=1.241874150e-23 wub1=1.063934483e-24 pub1=-2.122749420e-29 uc1=1.300133761e-11 luc1=4.321566231e-17 wuc1=8.984674179e-18 puc1=-1.792611501e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.28 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.5211602+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.028610852 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8962 eta0=0.08 etab=-0.07 u0=0.0309407 ua=-7.0410128e-10 ub=1.59378e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.396324 ags=0.4429907 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.29 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.169427526e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.353663987e-8 k1=5.483501070e-01 lk1=2.478842258e-8 k2=-2.468599297e-02 lk2=-3.121001191e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077667525e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.605073263e-8 nfactor=2.688232262e+00 lnfactor=1.653734701e-6 eta0=0.08 etab=-0.07 u0=3.131810464e-02 lu0=-3.001076750e-9 ua=-7.579478618e-10 lua=4.281816107e-16 ub=1.687370422e-18 lub=-7.442198968e-25 uc=8.117378080e-11 luc=-8.112334692e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.549110635e+00 la0=-1.214941142e-6 ags=4.327046453e-01 lags=8.179348265e-8 a1=0.0 a2=0.42385546 b0=4.189249708e-24 lb0=-1.655541632e-29 b1=0.0 keta=-1.056965338e-02 lketa=3.905767835e-8 dwg=0.0 dwb=0.0 pclm=-3.169121138e-01 lpclm=3.184275988e-06 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=1.446243820e-03 lpdiblc2=8.081444813e-9 pdiblcb=-4.968319824e+00 lpdiblcb=1.953541169e-5 drout=0.56 pscbe1=7.871095635e+08 lpscbe1=5.094147091e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141467060e-01 lkt1=-1.744081253e-8 kt2=-3.997479494e-02 lkt2=-8.642637524e-9 at=140000.0 ute=-1.817271588e+00 lute=2.144748568e-7 ua1=3.745936823e-10 lua1=-3.476059996e-16 ub1=-4.986867121e-19 lub1=5.846756647e-25 uc1=3.327652623e-12 luc1=9.414772148e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.30 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.174975316e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.134421944e-8 k1=5.404459826e-01 lk1=5.602458147e-8 k2=-2.491506218e-02 lk2=-3.030475765e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064178854e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.072017044e-8 nfactor=3.370399123e+00 lnfactor=-1.042107554e-6 eta0=0.08 etab=-0.07 u0=3.091862686e-02 lu0=-1.422388105e-9 ua=-5.069570504e-10 lua=-5.637042079e-16 ub=1.299150059e-18 lub=7.899807777e-25 uc=5.726534211e-11 luc=1.335995769e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=9.858058957e-01 la0=1.011172156e-6 ags=2.158259739e-01 lags=9.388721838e-7 a1=0.0 a2=0.42385546 b0=-2.056599416e-24 lb0=8.127436155e-30 b1=0.0 keta=-1.735957830e-03 lketa=4.147964760e-9 dwg=0.0 dwb=0.0 pclm=4.740059450e-01 lpclm=5.866193894e-8 pdiblc1=0.39 pdiblc2=2.166173716e-03 lpdiblc2=5.236367537e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.081380067e+08 lpscbe1=-3.216043418e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.150856518e-01 lkt1=-1.373021056e-8 kt2=-4.269599381e-02 lkt2=2.111216570e-9 at=1.643009184e+05 lat=-9.603433791e-2 ute=-1.936131845e+00 lute=6.841964476e-7 ua1=3.247381814e-11 lua1=1.004410991e-15 ub1=-2.950781812e-19 lub1=-2.199610200e-25 uc1=9.861007087e-12 luc1=6.832868211e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.31 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.979362322e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.952554794e-8 k1=6.287345350e-01 lk1=-1.163041665e-7 k2=-6.081372291e-02 lk2=3.976515613e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.965807302e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.103060895e-8 nfactor=3.356611396e+00 lnfactor=-1.015195551e-6 eta0=1.537410312e-01 leta0=-1.439337178e-7 etab=-5.631671063e-02 letab=-2.670815255e-8 u0=3.442203908e-02 lu0=-8.260631853e-9 ua=-1.431117554e-10 lua=-1.273886926e-15 ub=1.108883840e-18 lub=1.161357797e-24 uc=5.386395292e-11 luc=1.999906463e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.420255462e+04 lvsat=-8.202886504e-3 a0=2.036960762e+00 la0=-1.040557055e-6 ags=2.566041205e-01 lags=8.592780941e-7 a1=0.0 a2=0.42385546 b0=4.113198831e-24 lb0=-3.915275817e-30 b1=0.0 keta=4.960535517e-02 lketa=-9.606416860e-08 wketa=6.938893904e-24 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=1.374335140e-01 lpclm=7.156112720e-7 pdiblc1=1.705248073e-01 lpdiblc1=4.283894585e-7 pdiblc2=6.342319838e-03 lpdiblc2=-2.914972732e-9 pdiblcb=-4.861457464e-02 lpdiblcb=4.609283956e-8 drout=8.455643000e-01 ldrout=-5.573875314e-7 pscbe1=1.145718696e+09 lpscbe1=-6.910777669e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.585827200e-09 lalpha0=5.350920302e-14 alpha1=6.396342990e-01 lalpha1=4.106088148e-7 beta0=1.322319161e+01 lbeta0=1.242974195e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.860578468e-01 lkt1=1.247990683e-07 wkt1=4.440892099e-22 kt2=-4.711907459e-02 lkt2=1.074454392e-8 at=1.621895531e+05 lat=-9.191320394e-2 ute=-1.977870160e+00 lute=7.656646724e-7 ua1=-4.878066519e-10 lua1=2.019936555e-15 pua1=-8.271806126e-37 ub1=5.834418662e-19 lub1=-1.934727609e-24 uc1=1.020383967e-10 luc1=-1.115906132e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.32 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.732000160e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.116617845e-9 k1=4.427124355e-01 lk1=6.076673566e-8 k2=-2.190265573e-04 lk2=-1.791378402e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.968530194e-01 ldsub=6.010841108e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.286641533e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.863842250e-9 nfactor=1.882665198e+00 lnfactor=3.878258300e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-1.526556659e-22 peta0=-1.908195824e-28 etab=-1.600650675e-01 letab=7.204793714e-8 u0=2.861319205e-02 lu0=-2.731300735e-9 ua=-1.380653626e-09 lua=-9.589433327e-17 ub=2.406447592e-18 lub=-7.376848489e-26 wub=3.081487911e-39 uc=7.403259758e-11 luc=8.009149789e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.586375634e+04 lvsat=3.780989714e-2 a0=4.411313831e-01 la0=4.784826095e-7 ags=1.136653649e+00 lags=2.157566882e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.554655739e-02 lketa=1.354674908e-8 dwg=0.0 dwb=0.0 pclm=1.331358446e+00 lpclm=-4.208631858e-7 pdiblc1=7.295365653e-01 lpdiblc1=-1.037232127e-07 wpdiblc1=8.881784197e-22 pdiblc2=5.255966467e-03 lpdiblc2=-1.880893598e-9 pdiblcb=2.222914927e-02 lpdiblcb=-2.134195520e-08 wpdiblcb=-6.505213035e-24 ppdiblcb=3.469446952e-30 drout=-4.087838800e-01 ldrout=6.366026685e-7 pscbe1=7.601058167e+07 lpscbe1=3.271570623e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.816247674e-06 lalpha0=2.736703255e-12 walpha0=7.411538288e-28 palpha0=1.323488980e-33 alpha1=1.270731402e+00 lalpha1=-1.901205267e-7 beta0=1.137577438e+01 lbeta0=3.001495554e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.330485209e-01 lkt1=-2.084760183e-8 kt2=-3.484510072e-02 lkt2=-9.388186018e-10 at=8.283445085e+04 lat=-1.637658988e-2 ute=-1.101602841e+00 lute=-6.843753974e-8 ua1=2.169780508e-09 lua1=-5.097701682e-16 ub1=-2.235363667e-18 lub1=7.484398209e-25 uc1=-7.594942592e-11 luc1=5.783261332e-17 wuc1=2.584939414e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.33 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.125333257e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.989059316e-8 k1=4.142983009e-01 lk1=7.360654324e-8 k2=-5.123014741e-03 lk2=-1.569776494e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.331531951e-01 ldsub=8.889315138e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.348874771e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.051640481e-9 nfactor=2.604715256e+00 lnfactor=6.154512750e-8 eta0=0.49 etab=-0.000625 u0=2.667092004e-02 lu0=-1.853624917e-9 ua=-1.192661939e-09 lua=-1.808442046e-16 ub=2.017408214e-18 lub=1.020310179e-25 uc=7.692988093e-11 luc=-5.083123204e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.072438697e+05 lvsat=5.554580145e-3 a0=1.5 ags=2.125059674e+00 lags=-4.250662343e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.205412753e-02 lketa=-1.587843621e-9 dwg=0.0 dwb=0.0 pclm=4.635279131e-01 lpclm=-2.870705689e-8 pdiblc1=7.782704528e-01 lpdiblc1=-1.257451305e-07 wpdiblc1=-8.881784197e-22 pdiblc2=-1.078606283e-04 lpdiblc2=5.429179532e-10 pdiblcb=1.365048000e-01 lpdiblcb=-7.298095053e-08 wpdiblcb=5.551115123e-23 ppdiblcb=-2.775557562e-29 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.191548560e-06 lalpha0=2.189428516e-14 alpha1=0.85 beta0=1.712245588e+01 lbeta0=4.046793707e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.057206144e-01 lkt1=1.199153647e-8 kt2=-5.292091023e-02 lkt2=7.229296276e-09 wkt2=5.551115123e-23 at=6.589423514e+04 lat=-8.721628268e-3 ute=-2.038377412e+00 lute=3.548730904e-7 ua1=-4.578267072e-11 lua1=4.914007367e-16 ub1=1.195109989e-19 lub1=-3.156832979e-25 uc1=5.305567625e-11 luc1=-4.623412548e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.34 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.171028788e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.956310090e-08 wvth0=6.498750770e-07 pvth0=-1.311974304e-13 k1=5.374248511e-01 lk1=4.874963215e-8 k2=1.944997723e-02 lk2=-2.065858513e-08 wk2=-1.684127831e-07 pk2=3.399934107e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=7.898337811e-01 ldsub=-4.367818201e-08 wdsub=5.590371917e-11 pdsub=-1.128589873e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.170767983e-02 lcdscd=-1.273400711e-09 wcdscd=1.387778781e-23 cit=0.0 voff='-1.714711354e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.333905039e-09 wvoff=2.884586643e-07 pvoff=-5.823432360e-14 nfactor=6.184406878e+00 lnfactor=-6.611265968e-07 wnfactor=-6.739340461e-06 pnfactor=1.360544792e-12 eta0=1.411859226e+00 leta0=-1.861058623e-07 weta0=1.380618109e-14 peta0=-2.787205799e-21 etab=1.215937752e-01 letab=-2.467364857e-08 wetab=-8.106039279e-08 petab=1.636455316e-14 u0=-5.585034279e-03 lu0=4.658239396e-09 wu0=1.456099503e-08 pu0=-2.939588238e-15 ua=-3.791337613e-09 lua=3.437790392e-16 wua=-1.278882450e-16 pua=2.581820679e-23 ub=2.636456285e-18 lub=-2.294302563e-26 wub=1.563516123e-24 pub=-3.156441984e-31 uc=1.876506988e-10 luc=-2.286074176e-17 wuc=-2.568968277e-16 puc=5.186258847e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.878278900e+05 lvsat=-1.071380246e-02 wvsat=-1.499555026e-01 pvsat=3.027316681e-8 a0=1.5 ags=-2.298690174e+00 lags=4.680048089e-07 wags=-8.326672685e-22 pags=6.938893904e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.412227578e-01 lketa=-5.675725451e-08 wketa=-7.826181187e-07 pketa=1.579957284e-13 dwg=0.0 dwb=0.0 pclm=6.059181305e-02 lpclm=5.263808592e-08 wpclm=1.155758469e-06 ppclm=-2.333256755e-13 pdiblc1=-2.243565331e-01 lpdiblc1=7.666620805e-8 pdiblc2=-8.392336117e-03 lpdiblc2=2.215396149e-09 ppdiblc2=8.673617380e-31 pdiblcb=-4.542925080e-01 lpdiblcb=4.628980080e-8 drout=1.935739668e+00 ldrout=-1.889080599e-7 pscbe1=8.161650687e+08 lpscbe1=-3.263420225e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=9.460726714e-06 lalpha0=-1.243733670e-12 alpha1=0.85 beta0=2.684483517e+01 lbeta0=-1.558084282e-06 wbeta0=4.413451513e-06 pbeta0=-8.909920049e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.998761439e-01 lkt1=-9.376451085e-09 wkt1=-1.131654234e-07 pkt1=2.284594884e-14 kt2=5.059333590e-03 lkt2=-4.475813327e-9 at=-1.337710418e+05 lat=3.158699752e-02 wat=1.697481351e-01 pat=-3.426892327e-8 ute=1.676002233e+00 lute=-3.949895867e-7 ua1=6.932901369e-09 lua1=-9.174629760e-16 ub1=-5.498507054e-18 lub1=8.184878046e-25 uc1=-1.308925445e-10 luc1=3.667330950e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.35 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='1.375059692e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.067732016e-07 wvth0=-1.965247555e-06 pvth0=2.136875574e-13 k1=0.90707349 k2=-2.958942934e-01 lk2=2.092933262e-08 wk2=4.069974344e-07 pk2=-4.188633382e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586902379e-01 ldsub=-6.640391982e-12 wdsub=-1.304420114e-10 pdsub=1.328956256e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.310263022e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.531085334e-7 nfactor=-8.870386521e+00 lnfactor=1.324314611e-06 wnfactor=2.367387113e-05 pnfactor=-2.650379967e-12 eta0=6.941548766e-04 leta0=-1.639934862e-15 weta0=-3.221442386e-14 peta0=3.282037718e-21 etab=-6.549646949e-02 wetab=4.302535995e-8 u0=7.072192288e-02 lu0=-5.405198421e-09 wu0=-8.975373379e-08 pu0=1.081754251e-14 ua=-1.451891408e-09 lua=3.525053428e-17 wua=6.028150144e-16 pua=-7.054766976e-23 ub=6.970181767e-18 lub=-5.944790759e-25 wub=-9.851230895e-24 pub=1.189744053e-30 uc=1.430698928e-11 wuc=1.363560933e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.645626318e+03 lvsat=1.427415434e-02 wvsat=2.962069161e-01 pvsat=-2.856717912e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.940333415e-01 lketa=9.296145512e-08 wketa=1.826108944e-06 pketa=-1.860458053e-13 dwg=0.0 dwb=0.0 pclm=1.435665466e+00 lpclm=-1.287080025e-07 wpclm=-2.566626351e-06 ppclm=2.575861570e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.900562551e+01 lbeta0=-5.242414723e-07 wbeta0=-1.029805353e-05 pbeta0=1.049175992e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.709739600e-01 wkt1=6.006611748e-8 kt2=-0.028878939 at=2.586291603e+05 lat=-2.016313355e-02 wat=-3.960789819e-01 pat=4.035292276e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.36 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.166481222e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.002443909e-8 k1=5.401427619e-01 lk1=2.259480306e-7 k2=-2.486796516e-02 lk2=-7.467763289e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.036646356e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.157242546e-8 nfactor=2.875210105e+00 lnfactor=4.187878874e-7 eta0=0.08 etab=-0.07 u0=3.163311666e-02 lu0=-1.381501472e-8 ua=-7.265340304e-10 lua=4.475755662e-16 ub=1.636921731e-18 lub=-8.607586758e-25 uc=4.075029938e-11 luc=6.029797744e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.314757018e+00 la0=1.627414716e-6 ags=4.212090612e-01 lags=4.345846663e-7 a1=0.0 a2=0.42385546 b0=-5.255574854e-25 lb0=5.253045924e-29 b1=0.0 keta=-6.318895283e-03 lketa=1.318809922e-8 dwg=0.0 dwb=0.0 pclm=7.522374929e-02 lpclm=1.657452776e-7 pdiblc1=0.39 pdiblc2=3.376037021e-03 lpdiblc2=-1.822603774e-8 pdiblcb=5.951584812e-01 lpdiblcb=-6.198600671e-05 wpdiblcb=-2.775557562e-22 ppdiblcb=-2.042810365e-26 drout=0.56 pscbe1=6.698434685e+08 lpscbe1=2.467495241e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.264101520e-01 lkt1=2.009184746e-7 kt2=-4.661878793e-02 lkt2=1.108751152e-7 at=140000.0 ute=-1.906993821e+00 lute=2.328261231e-6 ua1=2.411981748e-10 lua1=1.789321105e-15 ub1=-5.159787779e-19 lub1=1.812005449e-24 uc1=1.749070723e-11 luc1=-4.635570604e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.37 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.5211602+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.028610852 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8962 eta0=0.08 etab=-0.07 u0=0.0309407 ua=-7.0410128e-10 ub=1.59378e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.396324 ags=0.4429907 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.38 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.169427526e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.353663987e-8 k1=5.483501070e-01 lk1=2.478842258e-8 k2=-2.468599297e-02 lk2=-3.121001191e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077667525e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.605073263e-8 nfactor=2.688232262e+00 lnfactor=1.653734701e-6 eta0=0.08 etab=-0.07 u0=3.131810464e-02 lu0=-3.001076750e-9 ua=-7.579478618e-10 lua=4.281816107e-16 ub=1.687370422e-18 lub=-7.442198968e-25 uc=8.117378080e-11 luc=-8.112334692e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.549110635e+00 la0=-1.214941142e-6 ags=4.327046453e-01 lags=8.179348265e-8 a1=0.0 a2=0.42385546 b0=4.189249708e-24 lb0=-1.655541632e-29 b1=0.0 keta=-1.056965338e-02 lketa=3.905767835e-8 dwg=0.0 dwb=0.0 pclm=-3.169121138e-01 lpclm=3.184275988e-06 wpclm=-2.220446049e-22 ppclm=-2.664535259e-27 pdiblc1=0.39 pdiblc2=1.446243820e-03 lpdiblc2=8.081444813e-9 pdiblcb=-4.968319824e+00 lpdiblcb=1.953541169e-5 drout=0.56 pscbe1=7.871095635e+08 lpscbe1=5.094147091e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141467060e-01 lkt1=-1.744081253e-8 kt2=-3.997479494e-02 lkt2=-8.642637524e-9 at=140000.0 ute=-1.817271588e+00 lute=2.144748568e-7 ua1=3.745936823e-10 lua1=-3.476059996e-16 wua1=-8.271806126e-31 ub1=-4.986867121e-19 lub1=5.846756647e-25 uc1=3.327652623e-12 luc1=9.414772148e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.39 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.174975316e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.134421944e-8 k1=5.404459826e-01 lk1=5.602458147e-8 k2=-2.491506218e-02 lk2=-3.030475765e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064178854e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.072017044e-8 nfactor=3.370399123e+00 lnfactor=-1.042107554e-6 eta0=0.08 etab=-0.07 u0=3.091862686e-02 lu0=-1.422388105e-9 ua=-5.069570504e-10 lua=-5.637042079e-16 ub=1.299150059e-18 lub=7.899807777e-25 uc=5.726534211e-11 luc=1.335995769e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=9.858058957e-01 la0=1.011172156e-6 ags=2.158259739e-01 lags=9.388721838e-7 a1=0.0 a2=0.42385546 b0=-2.056599416e-24 lb0=8.127436155e-30 b1=0.0 keta=-1.735957830e-03 lketa=4.147964760e-09 wketa=-1.734723476e-24 dwg=0.0 dwb=0.0 pclm=4.740059450e-01 lpclm=5.866193894e-8 pdiblc1=0.39 pdiblc2=2.166173716e-03 lpdiblc2=5.236367537e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.081380067e+08 lpscbe1=-3.216043418e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.150856518e-01 lkt1=-1.373021056e-8 kt2=-4.269599381e-02 lkt2=2.111216570e-9 at=1.643009184e+05 lat=-9.603433791e-2 ute=-1.936131845e+00 lute=6.841964476e-7 ua1=3.247381814e-11 lua1=1.004410991e-15 ub1=-2.950781812e-19 lub1=-2.199610200e-25 uc1=9.861007087e-12 luc1=6.832868211e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.40 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.979362322e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.952554794e-8 k1=6.287345350e-01 lk1=-1.163041665e-7 k2=-6.081372291e-02 lk2=3.976515613e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.965807302e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.103060895e-8 nfactor=3.356611396e+00 lnfactor=-1.015195551e-6 eta0=1.537410312e-01 leta0=-1.439337178e-7 etab=-5.631671062e-02 letab=-2.670815255e-8 u0=3.442203908e-02 lu0=-8.260631853e-9 ua=-1.431117554e-10 lua=-1.273886926e-15 ub=1.108883840e-18 lub=1.161357797e-24 uc=5.386395292e-11 luc=1.999906463e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.420255462e+04 lvsat=-8.202886504e-3 a0=2.036960762e+00 la0=-1.040557055e-6 ags=2.566041205e-01 lags=8.592780941e-7 a1=0.0 a2=0.42385546 b0=4.113198831e-24 lb0=-3.915275817e-30 b1=0.0 keta=4.960535517e-02 lketa=-9.606416860e-08 wketa=2.428612866e-23 pketa=1.101549407e-28 dwg=0.0 dwb=0.0 pclm=1.374335140e-01 lpclm=7.156112720e-7 pdiblc1=1.705248073e-01 lpdiblc1=4.283894585e-7 pdiblc2=6.342319838e-03 lpdiblc2=-2.914972732e-9 pdiblcb=-4.861457464e-02 lpdiblcb=4.609283956e-8 drout=8.455643000e-01 ldrout=-5.573875314e-7 pscbe1=1.145718696e+09 lpscbe1=-6.910777669e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.585827200e-09 lalpha0=5.350920302e-14 alpha1=6.396342990e-01 lalpha1=4.106088148e-7 beta0=1.322319161e+01 lbeta0=1.242974195e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.860578468e-01 lkt1=1.247990683e-7 kt2=-4.711907459e-02 lkt2=1.074454392e-8 at=1.621895531e+05 lat=-9.191320394e-2 ute=-1.977870160e+00 lute=7.656646724e-7 ua1=-4.878066519e-10 lua1=2.019936555e-15 pua1=-1.654361225e-36 ub1=5.834418662e-19 lub1=-1.934727609e-24 pub1=1.540743956e-45 uc1=1.020383967e-10 luc1=-1.115906132e-16 wuc1=-1.033975766e-31 puc1=-1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.41 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.732000160e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.116617845e-9 k1=4.427124355e-01 lk1=6.076673566e-8 k2=-2.190265573e-04 lk2=-1.791378402e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.968530194e-01 ldsub=6.010841108e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.286641533e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.863842250e-9 nfactor=1.882665198e+00 lnfactor=3.878258300e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-3.469446952e-22 peta0=2.116362641e-28 etab=-1.600650675e-01 letab=7.204793714e-8 u0=2.861319205e-02 lu0=-2.731300735e-9 ua=-1.380653626e-09 lua=-9.589433327e-17 ub=2.406447592e-18 lub=-7.376848489e-26 uc=7.403259758e-11 luc=8.009149789e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.586375634e+04 lvsat=3.780989714e-2 a0=4.411313831e-01 la0=4.784826095e-7 ags=1.136653649e+00 lags=2.157566882e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.554655739e-02 lketa=1.354674908e-8 dwg=0.0 dwb=0.0 pclm=1.331358446e+00 lpclm=-4.208631858e-7 pdiblc1=7.295365653e-01 lpdiblc1=-1.037232127e-7 pdiblc2=5.255966467e-03 lpdiblc2=-1.880893598e-9 pdiblcb=2.222914927e-02 lpdiblcb=-2.134195520e-08 wpdiblcb=-6.071532166e-24 ppdiblcb=-7.589415207e-30 drout=-4.087838800e-01 ldrout=6.366026685e-07 pdrout=-4.440892099e-28 pscbe1=7.601058167e+07 lpscbe1=3.271570623e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.816247674e-06 lalpha0=2.736703255e-12 walpha0=4.235164736e-28 alpha1=1.270731402e+00 lalpha1=-1.901205267e-7 beta0=1.137577438e+01 lbeta0=3.001495554e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.330485209e-01 lkt1=-2.084760183e-8 kt2=-3.484510072e-02 lkt2=-9.388186018e-10 at=8.283445085e+04 lat=-1.637658988e-2 ute=-1.101602841e+00 lute=-6.843753974e-8 ua1=2.169780508e-09 lua1=-5.097701682e-16 ub1=-2.235363667e-18 lub1=7.484398209e-25 uc1=-7.594942592e-11 luc1=5.783261332e-17 wuc1=5.169878828e-32 puc1=2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.42 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.125333257e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.989059316e-8 k1=4.142983009e-01 lk1=7.360654324e-8 k2=-5.123014741e-03 lk2=-1.569776494e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.331531951e-01 ldsub=8.889315138e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.348874771e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.051640481e-9 nfactor=2.604715256e+00 lnfactor=6.154512750e-8 eta0=0.49 etab=-0.000625 u0=2.667092004e-02 lu0=-1.853624917e-9 ua=-1.192661939e-09 lua=-1.808442046e-16 ub=2.017408214e-18 lub=1.020310179e-25 uc=7.692988093e-11 luc=-5.083123204e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.072438697e+05 lvsat=5.554580145e-3 a0=1.5 ags=2.125059674e+00 lags=-4.250662343e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.205412753e-02 lketa=-1.587843621e-9 dwg=0.0 dwb=0.0 pclm=4.635279131e-01 lpclm=-2.870705689e-8 pdiblc1=7.782704528e-01 lpdiblc1=-1.257451305e-7 pdiblc2=-1.078606283e-04 lpdiblc2=5.429179532e-10 pdiblcb=1.365048000e-01 lpdiblcb=-7.298095053e-8 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.191548560e-06 lalpha0=2.189428516e-14 alpha1=0.85 beta0=1.712245588e+01 lbeta0=4.046793707e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.057206144e-01 lkt1=1.199153647e-8 kt2=-5.292091023e-02 lkt2=7.229296276e-9 at=6.589423514e+04 lat=-8.721628268e-3 ute=-2.038377412e+00 lute=3.548730904e-7 ua1=-4.578267072e-11 lua1=4.914007367e-16 ub1=1.195109989e-19 lub1=-3.156832979e-25 uc1=5.305567625e-11 luc1=-4.623412548e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.43 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.918068443e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.589441037e-08 wvth0=1.001039874e-07 pvth0=-2.020909307e-14 k1=5.374248511e-01 lk1=4.874963215e-8 k2=-8.871542099e-02 lk2=1.177953628e-09 wk2=4.806100798e-08 pk2=-9.702604352e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=7.898617145e-01 ldsub=-4.368382123e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.170767983e-02 lcdscd=-1.273400711e-9 cit=0.0 voff='-2.733707583e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.376402303e-8 nfactor=1.965561723e+00 lnfactor=1.905780819e-07 wnfactor=1.703927162e-06 pnfactor=-3.439905195e-13 eta0=1.411859233e+00 leta0=-1.861058637e-7 etab=8.109035161e-02 letab=-1.649677690e-08 wetab=1.040834086e-23 petab=1.214306433e-29 u0=-4.451587590e-03 lu0=4.429418045e-09 wu0=1.229260324e-08 pu0=-2.481643034e-15 ua=-3.803319985e-09 lua=3.461980524e-16 wua=-1.039076615e-16 pua=2.097698262e-23 ub=2.574018250e-18 lub=-1.033797267e-26 wub=1.688474736e-24 pub=-3.408709682e-31 uc=-1.202484603e-10 luc=3.929824838e-17 wuc=3.593085333e-16 puc=-7.253756600e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.895465263e+05 lvsat=-1.106076249e-02 wvsat=-1.533950473e-01 pvsat=3.096754555e-8 a0=1.5 ags=-2.298690174e+00 lags=4.680048089e-07 wags=1.665334537e-21 pags=3.885780586e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.321449899e-01 lketa=5.899479977e-08 wketa=3.648753689e-07 pketa=-7.366140435e-14 dwg=0.0 dwb=0.0 pclm=5.167293187e-01 lpclm=-3.944740985e-08 wpclm=2.428804443e-07 ppclm=-4.903294697e-14 pdiblc1=-2.243565331e-01 lpdiblc1=7.666620805e-8 pdiblc2=-8.392336117e-03 lpdiblc2=2.215396149e-9 pdiblcb=-4.542925080e-01 lpdiblcb=4.628980080e-08 wpdiblcb=-8.881784197e-22 drout=1.935739668e+00 ldrout=-1.889080599e-7 pscbe1=8.161650687e+08 lpscbe1=-3.263420225e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=9.460726714e-06 lalpha0=-1.243733670e-12 alpha1=0.85 beta0=2.865414891e+01 lbeta0=-1.923350349e-06 wbeta0=7.924321184e-07 pbeta0=-1.599769885e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-5.844431246e-02 lkt1=-3.792885065e-08 wkt1=-3.962160592e-07 pkt1=7.998849424e-14 kt2=5.059333590e-03 lkt2=-4.475813327e-9 at=-4.895303898e+04 lat=1.446385428e-2 ute=1.676002233e+00 lute=-3.949895867e-07 wute=-1.776356839e-21 pute=2.220446049e-28 ua1=6.932901369e-09 lua1=-9.174629760e-16 ub1=-5.498507054e-18 lub1=8.184878046e-25 wub1=-6.162975822e-39 uc1=-1.308925445e-10 luc1=3.667330950e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.44 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.196341252e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=-5.313334836e-8 k1=0.90707349 k2=-7.978347759e-02 wk2=-2.550989573e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.410637829e+00 wnfactor=-9.044130798e-7 eta0=0.00069413878 etab=-0.043998 u0=2.913488844e-02 wu0=-6.524686850e-9 ua=-1.178240918e-09 wua=5.515226838e-17 ub=2.495629606e-18 wub=-8.962112172e-25 uc=1.777341785e-10 wuc=-1.907143359e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.056772617e+05 wvsat=8.141925912e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.151885894e-01 wketa=-1.936691094e-7 dwg=0.0 dwb=0.0 pclm=2.176156491e-01 wpclm=-1.289164557e-7 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.407016525e+01 wbeta0=-4.206083385e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.460433650e-01 wkt1=2.103041692e-7 kt2=-0.028878939 at=60720.487 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.45 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.073679991e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.644465785e-08 wvth0=1.560287507e-08 pvth0=2.630749350e-13 k1=4.477490672e-01 lk1=6.740104420e-06 wk1=1.553435516e-07 pk1=-1.095239445e-11 k2=7.805452917e-03 lk2=-2.441211891e-06 wk2=-5.493453662e-08 pk2=3.978906112e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016532196e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.579796916e-07 wvoff=-3.381838034e-09 pvoff=-5.036435645e-13 nfactor=2.656056846e+00 lnfactor=1.728070808e-05 wnfactor=3.684671955e-07 pnfactor=-2.835031738e-11 eta0=0.08 etab=-0.07 u0=3.272950912e-02 lu0=4.295285104e-08 wu0=-1.843388764e-09 pu0=-9.544506158e-14 ua=-7.630243481e-10 lua=-1.294657409e-15 wua=6.135197404e-17 pua=2.929254630e-21 ub=1.688423963e-18 lub=4.356375129e-24 wub=-8.659183710e-26 pub=-8.771681843e-30 uc=-8.384362722e-11 luc=5.795558838e-15 wuc=2.094825099e-16 puc=-8.730397417e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.038470972e+00 la0=9.646109697e-06 wa0=4.645258072e-07 pa0=-1.348200828e-11 ags=2.836420188e-01 lags=8.951591162e-06 wags=2.312944947e-07 pags=-1.431983040e-11 a1=0.0 a2=0.42385546 b0=-1.001074388e-23 lb0=3.680439064e-28 wb0=1.594765257e-29 pb0=-5.304797000e-34 b1=0.0 keta=-5.214759735e-03 lketa=-2.559776383e-07 wketa=-1.856407387e-09 pketa=4.525542762e-13 dwg=0.0 dwb=0.0 pclm=5.027584910e-02 lpclm=6.635028134e-07 wpclm=4.194545344e-08 ppclm=-8.368906956e-13 pdiblc1=0.39 pdiblc2=6.634586870e-03 lpdiblc2=-1.244542634e-07 wpdiblc2=-5.478671549e-09 ppdiblc2=1.786038528e-13 pdiblcb=1.014476295e+01 lpdiblcb=-2.700786015e-04 wpdiblcb=-1.605596009e-05 ppdiblcb=3.498706576e-10 drout=0.56 pscbe1=2.744684002e+08 lpscbe1=1.227348040e+04 wpscbe1=6.647528006e+02 ppscbe1=-1.648701858e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.387816291e-01 lkt1=-9.819013578e-07 wkt1=2.080043668e-08 pkt1=1.988701006e-12 kt2=-4.800972373e-02 lkt2=-1.085207796e-06 wkt2=2.338610957e-09 pkt2=2.011000512e-12 at=140000.0 ute=-1.881004968e+00 lute=-2.830527519e-05 wute=-4.369563036e-08 pute=5.150483872e-11 ua1=7.378678020e-10 lua1=-6.939996316e-14 wua1=-8.350615709e-16 pua1=1.196921098e-19 ub1=-1.175869020e-18 lub1=4.594990070e-23 wub1=1.109487982e-24 pub1=-7.421001432e-29 uc1=-5.173249802e-12 luc1=2.777144532e-15 wuc1=3.810540956e-17 puc1=-4.747213068e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.46 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.040377539e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.878834541e-8 k1=7.855670614e-01 wk1=-3.935968941e-7 k2=-1.145495216e-01 wk2=1.444905758e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.872312583e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-2.862474944e-8 nfactor=3.522176090e+00 wnfactor=-1.052467371e-6 eta0=0.08 etab=-0.07 u0=3.488233125e-02 wu0=-6.627151337e-9 ua=-8.279133382e-10 wua=2.081679374e-16 ub=1.906768045e-18 wub=-5.262336856e-25 uc=2.066331874e-10 wuc=-2.280901389e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.521939659e+00 wa0=-2.112003704e-7 ags=7.323010281e-01 wags=-4.864238194e-7 a1=0.0 a2=0.42385546 b0=8.435832978e-24 wb0=-1.064030172e-29 b1=0.0 keta=-1.804450939e-02 wketa=2.082587887e-8 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=3.968660562e-04 wpdiblc2=3.473058507e-9 pdiblcb=-3.391735258e+00 wpdiblcb=1.479762863e-6 drout=0.56 pscbe1=8.896224500e+08 wpscbe1=-1.615862587e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.879951022e-01 wkt1=1.204752997e-7 kt2=-1.024009761e-01 wkt2=1.031311383e-7 at=140000.0 ute=-3.299681993e+00 wute=2.537757152e-6 ua1=-2.740499133e-09 wua1=5.163977307e-15 ub1=1.127167004e-18 wub1=-2.609961543e-24 uc1=1.340188661e-10 wuc1=-1.998276990e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.47 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.906863338e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.061689032e-07 wvth0=4.414549452e-08 pvth0=-1.221182223e-13 k1=8.227477715e-01 lk1=-2.956565825e-07 wk1=-4.613508302e-07 pk1=5.387712368e-13 k2=-1.228611414e-01 lk2=6.609301178e-08 wk2=1.650640369e-07 pk2=-1.635977144e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.076022498e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.332003996e-08 wvoff=-4.540666885e-08 pvoff=1.334478261e-13 nfactor=3.170129836e+00 lnfactor=2.799429913e-06 wnfactor=-8.102249930e-07 pnfactor=-1.926282564e-12 eta0=0.08 etab=-0.07 u0=3.377999375e-02 lu0=8.765656625e-09 wu0=-4.139228329e-09 pu0=-1.978366769e-14 ua=-1.153238795e-09 lua=2.586949319e-15 wua=6.646113425e-16 pua=-3.629583641e-21 ub=2.293025369e-18 lub=-3.071472278e-24 wub=-1.018300987e-24 pub=3.912860628e-30 uc=2.462203393e-10 luc=-3.147923208e-16 wuc=-2.774964098e-16 puc=3.928727865e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.743644246e+00 la0=-1.762968497e-06 wa0=-3.270736397e-07 pa0=9.214104489e-13 ags=6.713011755e-01 lags=4.850635691e-07 wags=-4.011575952e-07 pags=-6.780268683e-13 a1=0.0 a2=0.42385546 b0=1.677018499e-23 lb0=-6.627377544e-29 wb0=-2.115260328e-29 pb0=8.359257099e-35 b1=0.0 keta=-4.199145147e-03 lketa=-1.100966888e-07 wketa=-1.071087564e-08 pketa=2.507765190e-13 dwg=0.0 dwb=0.0 pclm=-1.854434352e-01 lpclm=2.138852701e-06 wpclm=-2.210411815e-07 ppclm=1.757693172e-12 pdiblc1=0.39 pdiblc2=-3.095106662e-03 lpdiblc2=2.776775151e-08 wpdiblc2=7.635472475e-09 ppdiblc2=-3.309902055e-14 pdiblcb=-6.717969533e+00 lpdiblcb=2.644981913e-05 wpdiblcb=2.941724548e-06 ppdiblcb=-1.162534535e-11 drout=0.56 pscbe1=8.156586009e+08 lpscbe1=5.881517268e+02 wpscbe1=-4.800012455e+01 ppscbe1=-9.032234219e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.828644579e-01 lkt1=-4.079827256e-08 wkt1=1.155366680e-07 pkt1=3.927141142e-14 kt2=-9.823322323e-02 lkt2=-3.314147518e-08 wkt2=9.795117718e-08 pkt2=4.119043472e-14 at=140000.0 ute=-2.807721695e+00 lute=-3.912009749e-06 wute=1.665265555e-06 pute=6.937949350e-12 ua1=-2.263167420e-09 lua1=-3.795684975e-15 wua1=4.434925773e-15 pua1=5.797331040e-21 ub1=8.144035246e-19 lub1=2.487057972e-24 wub1=-2.207727503e-24 pub1=-3.198517225e-30 uc1=1.047914674e-10 luc1=2.324127960e-16 wuc1=-1.705933441e-16 puc1=-2.324681116e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.48 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.432798274e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.016743247e-07 wvth0=-4.334834119e-08 pvth0=2.236470047e-13 k1=8.352913552e-01 lk1=-3.452273326e-07 wk1=-4.957300116e-07 pk1=6.746336707e-13 k2=-1.447850732e-01 lk2=1.527337813e-07 wk2=2.015400867e-07 pk2=-3.077467224e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.657853173e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.726890067e-07 wvoff=9.981576925e-08 pvoff=-4.404539678e-13 nfactor=3.681868463e+00 lnfactor=7.770997557e-07 wnfactor=-5.236802542e-07 pnfactor=-3.058673273e-12 eta0=0.08 etab=-0.07 u0=3.465036219e-02 lu0=5.326064105e-09 wu0=-6.274248722e-09 pu0=-1.134632117e-14 ua=-1.272480459e-09 lua=3.058178187e-15 wua=1.287091349e-15 pua=-6.089550551e-21 ub=2.408638467e-18 lub=-3.528361483e-24 wub=-1.865407269e-24 pub=7.260523846e-30 uc=2.371972062e-10 luc=-2.791339728e-16 wuc=-3.025234017e-16 puc=4.917764802e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=-1.583371006e-01 la0=5.753435450e-06 wa0=1.923672791e-06 pa0=-7.973271606e-12 ags=2.351956722e-01 lags=2.208500622e-06 wags=-3.256669991e-08 pags=-2.134654224e-12 a1=0.0 a2=0.42385546 b0=-8.232871054e-24 lb0=3.253532669e-29 wb0=1.038430138e-29 pb0=-4.103752334e-35 b1=0.0 keta=-9.078413925e-02 lketa=2.320769042e-07 wketa=1.497186665e-07 pketa=-3.832219404e-13 dwg=0.0 dwb=0.0 pclm=3.664938643e-01 lpclm=-4.233782640e-08 wpclm=1.807624265e-07 ppclm=1.698131275e-13 pdiblc1=0.39 pdiblc2=4.348969113e-03 lpdiblc2=-1.650350109e-09 wpdiblc2=-3.669981923e-09 ppdiblc2=1.157878989e-14 pdiblcb=-0.025 drout=0.56 pscbe1=1.157593969e+09 lpscbe1=-7.631361590e+02 wpscbe1=-5.875479980e+02 ppscbe1=1.229005568e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.733301761e-01 lkt1=-7.847661976e-08 wkt1=9.792780007e-08 pkt1=1.088595622e-13 kt2=-9.996658525e-02 lkt2=-2.629143476e-08 wkt2=9.629030535e-08 pkt2=4.775400253e-14 at=1.528704342e+05 lat=-5.086242451e-02 wat=1.921832458e-02 pat=-7.594853178e-8 ute=-2.547434600e+00 lute=-4.940633374e-06 wute=1.027796771e-06 pute=9.457150125e-12 ua1=2.075577560e-09 lua1=-2.094188883e-14 wua1=-3.435115270e-15 pua1=3.689879670e-20 ub1=-3.573678942e-18 lub1=1.982823770e-23 wub1=5.512383589e-24 pub1=-3.370747757e-29 uc1=5.940793136e-11 luc1=4.117631299e-16 wuc1=-8.330433381e-17 puc1=-5.774238927e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.49 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.255010315e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.282158692e-07 wvth0=1.217868965e-07 pvth0=-9.867732824e-14 k1=7.249917915e-01 lk1=-1.299357099e-07 wk1=-1.618394430e-07 pk1=2.291901381e-14 k2=-9.347853572e-02 lk2=5.258952558e-08 wk2=5.492006841e-08 pk2=-2.156189448e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.621737396e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.020773982e-07 wvoff=-1.611974983e-07 pvoff=6.901286980e-14 nfactor=4.905492361e+00 lnfactor=-1.611268481e-06 wnfactor=-2.604167642e-06 pnfactor=1.002190530e-12 eta0=1.537411742e-01 leta0=-1.439339967e-07 weta0=-2.403146453e-13 peta0=4.690655904e-19 etab=-5.631671062e-02 letab=-2.670815255e-8 u0=4.915098778e-02 lu0=-2.297743146e-08 wu0=-2.476410549e-08 pu0=2.474367896e-14 ua=2.233013691e-09 lua=-3.784129240e-15 wua=-3.995031987e-15 pua=4.220525628e-21 ub=-1.432272381e-18 lub=3.968639423e-24 wub=4.272501859e-24 pub=-4.719944359e-30 uc=9.905424606e-11 luc=-9.495353580e-18 wuc=-7.597943405e-17 puc=4.958961421e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.254098381e+05 lvsat=-8.863460018e-02 wvsat=-6.928271226e-02 pvsat=1.352316097e-7 a0=3.909768631e+00 la0=-2.187022834e-06 wa0=-3.148793073e-06 pa0=1.927578137e-12 ags=1.103361330e-01 lags=2.452211584e-06 wags=2.459235853e-07 pags=-2.678234121e-12 a1=0.0 a2=0.42385546 b0=1.646574211e-23 lb0=-1.567342706e-29 wb0=-2.076860277e-29 pb0=1.976923837e-35 b1=0.0 keta=2.776841838e-01 lketa=-4.871294146e-07 wketa=-3.834739523e-07 pketa=6.575066016e-13 dwg=0.0 dwb=0.0 pclm=-7.477462322e-01 lpclm=2.132526247e-06 wpclm=1.488272181e-06 ppclm=-2.382290320e-12 pdiblc1=-6.352265768e-01 lpdiblc1=2.001120276e-06 wpdiblc1=1.354727529e-06 ppdiblc1=-2.644266924e-12 pdiblc2=1.093904860e-02 lpdiblc2=-1.451340105e-08 wpdiblc2=-7.728581195e-09 ppdiblc2=1.950069269e-14 pdiblcb=-1.892049255e-01 lpdiblcb=3.205084741e-07 wpdiblcb=2.363776499e-07 ppdiblcb=-4.613810436e-13 drout=1.238054913e+00 ldrout=-1.323482502e-06 wdrout=-6.599031030e-07 pdrout=1.288052329e-12 pscbe1=2.183962974e+09 lpscbe1=-2.766486317e+03 wpscbe1=-1.745622946e+03 ppscbe1=3.489430055e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.317334756e-08 lalpha0=2.209009068e-13 walpha0=1.441887872e-13 palpha0=-2.814393542e-19 alpha1=-4.294967464e-01 lalpha1=2.497425389e-06 walpha1=1.797553547e-06 palpha1=-3.508610616e-12 beta0=1.131076201e+01 lbeta0=4.975809190e-06 wbeta0=3.215409955e-06 pbeta0=-6.276097599e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-5.693217365e-01 lkt1=3.040755831e-07 wkt1=3.081256095e-07 pkt1=-3.014215484e-13 kt2=-1.884375369e-01 lkt2=1.463933349e-07 wkt2=2.376018397e-07 pkt2=-2.280692965e-13 at=2.424662890e+05 lat=-2.257428711e-01 wat=-1.349710422e-01 pat=2.250107637e-7 ute=-8.433700634e+00 lute=6.548657458e-06 wute=1.085432980e-05 pute=-9.723072996e-12 ua1=-1.955519357e-08 lua1=2.127880236e-14 wua1=3.205841711e-14 pua1=-3.238035477e-20 ub1=1.617999044e-17 lub1=-1.872857426e-23 wub1=-2.622282025e-23 pub1=2.823586383e-29 uc1=6.372039961e-10 luc1=-7.160260307e-16 wuc1=-8.997856959e-16 puc1=1.016250565e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.50 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.561446423e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.858698228e-09 wvth0=2.867557498e-08 pvth0=-1.004643037e-14 k1=5.615189451e-01 lk1=2.567098662e-08 wk1=-1.997519984e-07 pk1=5.900725497e-14 k2=-2.268402434e-02 lk2=-1.479842471e-08 wk2=3.777089500e-08 pk2=-5.237922152e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.520285266e-01 ldsub=1.027759941e-07 wdsub=7.536440578e-08 pdsub=-7.173794593e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.455146000e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.471388977e-08 wvoff=-1.414205217e-07 pvoff=5.018754159e-14 nfactor=4.836077604e+00 lnfactor=-1.545193893e-06 wnfactor=-4.965637255e-06 pnfactor=3.250028587e-12 eta0=-4.380247683e-01 leta0=4.193567603e-07 weta0=4.806292907e-13 peta0=-2.171872447e-19 etab=-1.592169017e-01 letab=7.124058419e-08 wetab=-1.426039892e-09 petab=1.357420278e-15 u0=2.703625902e-02 lu0=-1.926841337e-09 wu0=2.651332194e-09 pu0=-1.352555284e-15 ua=-1.583136910e-09 lua=-1.516079907e-16 wua=3.404396003e-16 pua=9.367259795e-23 ub=2.664920372e-18 lub=6.859948861e-26 wub=-4.345759726e-25 pub=-2.393664060e-31 uc=1.057843408e-10 luc=-1.590160287e-17 wuc=-5.338490439e-17 puc=2.808231072e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.111483594e+04 lvsat=8.891469306e-02 wvsat=1.630522407e-01 pvsat=-8.592361769e-8 a0=1.713580280e+00 la0=-9.651287052e-08 wa0=-2.139396324e-06 pa0=9.667525504e-13 ags=3.801960734e+00 lags=-1.061775733e-06 wags=-4.481239438e-06 pags=1.821462545e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.028197102e-01 lketa=1.606293125e-07 wketa=5.670647718e-07 pketa=-2.472931496e-13 dwg=0.0 dwb=0.0 pclm=2.751429902e+00 lpclm=-1.198273031e-06 wpclm=-2.387597382e-06 ppclm=1.307076275e-12 pdiblc1=1.369703661e+00 lpdiblc1=9.266527642e-08 wpdiblc1=-1.076327021e-06 ppdiblc1=-3.301922872e-13 pdiblc2=-7.799595524e-03 lpdiblc2=3.323558260e-09 wpdiblc2=2.195060360e-08 ppdiblc2=-8.750359408e-15 pdiblcb=3.034098510e-01 lpdiblcb=-1.484021719e-07 wpdiblcb=-4.727552997e-07 ppdiblcb=2.136291376e-13 drout=-1.193765107e+00 ldrout=9.913207702e-07 wdrout=1.319806206e-06 pdrout=-5.963953482e-13 pscbe1=-2.098236516e+09 lpscbe1=1.309658015e+03 wpscbe1=3.655609479e+03 ppscbe1=-1.651900467e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.135708887e-05 lalpha0=1.095232689e-11 walpha0=1.435990420e-11 palpha0=-1.381310875e-17 alpha1=3.408993493e+00 lalpha1=-1.156360539e-06 walpha1=-3.595107095e-06 palpha1=1.624560589e-12 beta0=3.915278132e+00 lbeta0=1.201542978e-05 wbeta0=1.254349648e-05 pbeta0=-1.515532592e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.005301102e-01 lkt1=-4.697015890e-08 wkt1=-5.467391924e-08 pkt1=4.392042990e-14 kt2=-3.103052505e-02 lkt2=-3.439408999e-09 wkt2=-6.413529991e-09 pkt2=4.204297649e-15 at=-2.239755128e+04 lat=2.637598604e-02 wat=1.769288803e-01 pat=-7.188084645e-8 ute=-1.752407620e+00 lute=1.888615829e-07 wute=1.094212393e-06 pute=-4.326026755e-13 ua1=4.528719309e-09 lua1=-1.646216717e-15 wua1=-3.966135703e-15 pua1=1.910732584e-21 ub1=-6.404124217e-18 lub1=2.768815392e-24 wub1=7.009028826e-24 pub1=-3.396901895e-30 uc1=-3.008165365e-10 luc1=1.768578919e-16 wuc1=3.780740201e-16 puc1=-2.001198195e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.51 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.845226536e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-8.964785863e-09 wvth0=4.709495931e-08 pvth0=-1.836980018e-14 k1=7.994915626e-01 lk1=-8.186431772e-08 wk1=-6.476339052e-07 pk1=2.613965789e-13 k2=-1.534059664e-01 lk2=4.427233717e-08 wk2=2.493113888e-07 pk2=-1.008290520e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-5.571655909e-02 ldsub=1.966520511e-07 wdsub=3.175508728e-07 pdsub=-1.811774088e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-2.719280928e-03 lcdscd=3.668948785e-09 wcdscd=1.365112565e-08 pcdscd=-6.168684310e-15 cit=0.0 voff='-1.833232664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.799445287e-08 wvoff=8.143615818e-08 pvoff=-5.051715777e-14 nfactor=-5.727328209e-01 lnfactor=8.989447709e-07 wnfactor=5.342313356e-06 pnfactor=-1.407938443e-12 eta0=-6.966223827e-01 leta0=5.362121089e-07 weta0=1.995094318e-06 peta0=-9.015452154e-13 etab=-1.075057916e-01 letab=4.787331606e-08 wetab=1.797010263e-07 petab=-8.049045950e-14 u0=5.476874060e-02 lu0=-1.445862284e-08 wu0=-4.724148386e-08 pu0=2.119306032e-14 ua=4.371757035e-10 lua=-1.064548875e-15 wua=-2.740281885e-15 pua=1.485792103e-21 ub=2.182538473e-18 lub=2.865787034e-25 wub=-2.776371374e-25 pub=-3.102840838e-31 uc=1.115228123e-10 luc=-1.849470910e-17 wuc=-5.816185647e-17 puc=3.024092460e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.647651524e+05 lvsat=-1.315618197e-02 wvsat=-9.671179819e-02 pvsat=3.145881598e-8 a0=1.5 ags=5.593287916e+00 lags=-1.871242451e-06 wags=-5.831208444e-06 pags=2.431487889e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.581875311e-01 lketa=5.008467877e-08 wketa=2.120708664e-07 pketa=-8.687814868e-14 dwg=0.0 dwb=0.0 pclm=-2.800006429e-01 lpclm=1.715728356e-07 wpclm=1.250110919e-06 ppclm=-3.367349894e-13 pdiblc1=3.209770237e+00 lpdiblc1=-7.388258479e-07 wpdiblc1=-4.088134079e-06 ppdiblc1=1.030786098e-12 pdiblc2=1.123720671e-02 lpdiblc2=-5.278810970e-09 wpdiblc2=-1.907471131e-08 ppdiblc2=9.788200916e-15 pdiblcb=4.316514050e-01 lpdiblcb=-2.063520935e-07 wpdiblcb=-4.962364802e-07 ppdiblcb=2.242398369e-13 drout=-2.044893600e-01 ldrout=5.442858565e-07 wdrout=2.025134460e-06 pdrout=-9.151197848e-13 pscbe1=7.791922328e+08 lpscbe1=9.402634663e+00 wpscbe1=3.498455681e+01 ppscbe1=-1.580885652e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.266577463e-05 lalpha0=9.685130335e-14 walpha0=-1.592922473e-11 palpha0=-1.260268837e-19 alpha1=0.85 beta0=2.803564484e+01 lbeta0=1.115894353e-06 wbeta0=-1.834858469e-05 pbeta0=-1.195781397e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.384323881e-01 lkt1=1.534526031e-08 wkt1=5.499902469e-08 pkt1=-5.638689673e-15 kt2=-8.456639466e-02 lkt2=2.075243329e-08 wkt2=5.320624917e-08 pkt2=-2.273674778e-14 at=6.131394926e+04 lat=-1.145165054e-02 wat=7.700935418e-03 pat=4.590046506e-9 ute=-4.704003976e+00 lute=1.522631896e-06 wute=4.481776586e-06 pute=-1.963378570e-12 ua1=-6.177530495e-09 lua1=3.191734151e-15 wua1=1.030944251e-14 pua1=-4.540129977e-21 ub1=5.884606908e-18 lub1=-2.784228718e-24 wub1=-9.692982584e-24 pub1=4.150419723e-30 uc1=3.565353589e-10 luc1=-1.201869399e-16 wuc1=-5.102470671e-16 puc1=2.012956017e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.52 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='8.584319749e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.426187355e-08 wvth0=-1.800465104e-07 pvth0=2.748574687e-14 k1=-5.726845787e-01 lk1=1.951519739e-07 wk1=1.866451407e-06 pk1=-2.461494780e-13 k2=4.068947626e-01 lk2=-6.884173429e-08 wk2=-7.852192971e-07 pk2=1.080230374e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.784571499e+00 ldsub=-1.748671423e-07 wdsub=-1.672427444e-06 pdsub=2.205614038e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=4.070511172e-02 lcdscd=-5.097611026e-09 wcdscd=-4.875402018e-08 pcdscd=6.429728935e-15 cit=0.0 voff='2.622033209e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.194890009e-08 wvoff=-4.868106389e-07 pvoff=6.420107387e-14 nfactor=5.585002960e+00 lnfactor=-3.441850863e-07 wnfactor=-4.381519016e-06 pnfactor=5.551185599e-13 eta0=5.649796314e+00 leta0=-7.450092439e-07 weta0=-7.125336849e-06 peta0=9.396965490e-13 etab=4.567491369e-01 letab=-6.603903317e-08 wetab=-6.316033803e-07 petab=8.329648539e-14 u0=-1.013327432e-01 lu0=1.705530081e-08 wu0=1.751810216e-07 pu0=-2.370981749e-14 ua=-1.173418409e-08 lua=1.392617413e-15 wua=1.323042865e-14 pua=-1.738390909e-21 ub=6.904551078e-18 lub=-6.667059232e-25 wub=-5.592545380e-24 pub=7.626949072e-31 uc=3.087113398e-11 luc=-2.212667638e-18 wuc=1.052278348e-16 puc=-2.744349656e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.315110571e+04 lvsat=2.881816014e-02 wvsat=2.378446008e-01 pvsat=-3.608176440e-8 a0=1.5 ags=-1.295593062e+01 lags=1.873492336e-06 wags=1.791825282e-05 pags=-2.363077101e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.592803113e-01 lketa=-3.419414674e-08 wketa=-6.295010015e-07 pketa=8.301922158e-14 dwg=0.0 dwb=0.0 pclm=1.377981681e+00 lpclm=-1.631422939e-07 wpclm=-1.205162100e-06 ppclm=1.589379829e-13 pdiblc1=-1.970172384e+00 lpdiblc1=3.069061482e-07 wpdiblc1=2.935278597e-06 ppdiblc1=-3.871074767e-13 pdiblc2=-5.884055588e-02 lpdiblc2=8.868557820e-09 wpdiblc2=8.481970175e-08 ppdiblc2=-1.118610709e-14 pdiblcb=-1.508387526e+00 lpdiblcb=1.853049059e-07 wpdiblcb=1.772273144e-06 ppdiblcb=-2.337291545e-13 drout=6.237487382e+00 ldrout=-7.562268502e-07 wdrout=-7.232623070e-06 pdrout=9.538455631e-13 pscbe1=8.904785230e+08 lpscbe1=-1.306395290e+01 wpscbe1=-1.249448458e+02 ppscbe1=1.647785120e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.785534461e-05 lalpha0=-4.988444272e-12 walpha0=-4.774049574e-11 palpha0=6.296064319e-18 alpha1=0.85 beta0=7.092920990e+01 lbeta0=-7.543501454e-06 wbeta0=-7.028555798e-05 pbeta0=9.289306708e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.405326468e-01 lkt1=1.576926264e-08 wkt1=7.806526330e-08 pkt1=-1.029532499e-14 kt2=1.069809761e-01 lkt2=-1.791734147e-08 wkt2=-1.713630999e-07 pkt2=2.259953697e-14 at=-2.143224274e+05 lat=4.419409682e-02 wat=2.780391909e-01 pat=-4.998611084e-8 ute=1.067056579e+01 lute=-1.581201624e-06 wute=-1.512275759e-05 pute=1.994404394e-12 ua1=2.782504468e-08 lua1=-3.672739728e-15 wua1=-3.512642018e-14 pua1=4.632507419e-21 ub1=-2.413682267e-17 lub1=3.276527506e-24 wub1=3.133701008e-23 pub1=-4.132756227e-30 uc1=-9.660042140e-10 luc1=1.468086716e-16 wuc1=1.404091622e-15 puc1=-1.851730073e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.53 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='3.711603167e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.836673235e-8 k1=0.90707349 k2=-1.151041174e-01 wk2=3.387547300e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.975187397e+00 wnfactor=-1.722806885e-7 eta0=0.00069413878 etab=-0.043998 u0=2.799066811e-02 wu0=-4.600884036e-9 ua=-1.174532494e-09 wua=4.891721307e-17 ub=1.849191146e-18 wub=1.906599882e-25 uc=1.409337496e-11 wuc=8.441854720e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.753652851e+05 wvsat=-3.574874778e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=0.0 dwg=0.0 dwb=0.0 pclm=0.14094 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.372990557e+01 wbeta0=1.514777448e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=1.207834394e+05 wat=-1.009851632e-1 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.54 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.590239303e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.636885092e-06 wvth0=-1.756840874e-07 pvth0=3.505228005e-12 k1=4.913208483e-01 lk1=-3.552406136e-07 wk1=1.003855055e-07 pk1=-2.002879660e-12 k2=1.758888301e-02 lk2=-3.508246201e-07 wk2=-6.727459224e-08 pk2=1.342254659e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.216279298e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.841650295e-07 wvoff=-1.535232189e-08 pvoff=3.063076993e-13 nfactor=3.013624176e+00 lnfactor=-6.501603257e-06 wnfactor=-8.254034387e-08 pnfactor=1.646835119e-12 eta0=0.08 etab=-0.07 u0=5.190747709e-02 lu0=-4.445134854e-07 wu0=-2.603298169e-08 pu0=5.194069528e-13 ua=9.853359250e-10 lua=-3.288488529e-14 wua=-2.143893302e-15 pua=4.277470405e-20 ub=6.132927897e-19 lub=1.748317910e-23 wub=1.269494765e-24 pub=-2.532880849e-29 uc=1.901892776e-10 luc=-3.279895256e-15 wuc=-1.361612217e-16 puc=2.716672492e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.569026678e+00 la0=-4.280290551e-06 wa0=-2.046757762e-07 pa0=4.083666731e-12 ags=9.390990363e-01 lags=-1.182037291e-05 wags=-5.954478614e-07 pags=1.188030487e-11 a1=0.0 a2=0.42385546 b0=-3.053957932e-07 lb0=6.093220525e-12 wb0=3.852024327e-13 pb0=-7.685513099e-18 b1=-1.212267661e-08 lb1=2.418702010e-13 wb1=1.529059870e-14 pb1=-3.050762057e-19 keta=-1.203383205e-02 lketa=2.095042146e-07 wketa=6.744638540e-09 pketa=-1.345682255e-13 dwg=0.0 dwb=0.0 pclm=4.042617819e-01 lpclm=-6.399182393e-06 wpclm=-4.045447913e-07 ppclm=8.071429534e-12 pdiblc1=0.39 pdiblc2=9.519222739e-03 lpdiblc2=-1.270705381e-07 wpdiblc2=-9.117126232e-09 ppdiblc2=1.819038176e-13 pdiblcb=-1.454963836e+01 lpdiblcb=2.460283836e-04 wpdiblcb=1.509163156e-05 ppdiblcb=-3.011064370e-10 drout=0.56 pscbe1=3.537042373e+09 lpscbe1=-5.537701580e+04 wpscbe1=-3.450403528e+03 ppscbe1=6.884204059e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.664501274e-01 lkt1=3.471031279e-06 wkt1=1.818315222e-07 pkt1=-3.627880894e-12 kt2=-1.017009639e-01 lkt2=1.617385465e-06 wkt2=7.006055340e-08 pkt2=-1.397839824e-12 at=-2.841060618e+04 lat=3.360108374e+00 wat=2.124200026e-01 pat=-4.238178614e-6 ute=-5.163085353e+00 lute=7.732122739e-05 wute=4.096064565e-06 pute=-8.172419276e-11 ua1=-3.726030223e-09 lua1=1.013481777e-13 wua1=4.795351213e-15 pua1=-9.567627676e-20 ub1=3.981350790e-19 lub1=-2.673941273e-23 wub1=-8.758380165e-25 pub1=1.747461588e-29 uc1=-6.470630903e-11 luc1=8.040206218e-16 wuc1=1.131957669e-16 puc1=-2.258468471e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.55 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.5268617+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.47351598 k2=5.34690000000056e-6 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.11141737+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.68776 eta0=0.08 etab=-0.07 u0=0.0296282 ua=-6.6287385e-10 ub=1.48956e-18 uc=2.5799e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.354496 ags=0.346655 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.0015333577 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0031503727 pdiblcb=-2.2185512 drout=0.56 pscbe1=761513800.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.29248 kt2=-0.020636654 at=140000.0 ute=-1.2877 ua1=1.3536e-9 ub1=-9.4206e-19 uc1=-2.4408323e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.56 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.256857190e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.351260879e-9 k1=4.569800848e-01 lk1=1.314914708e-7 k2=8.004757165e-03 lk2=-6.361035850e-08 wk2=1.877025011e-24 pk2=-2.442165394e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.167594931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.247992715e-8 nfactor=2.527768098e+00 lnfactor=1.272236568e-6 eta0=0.08 etab=-0.07 u0=3.049833504e-02 lu0=-6.919210278e-9 ua=-6.263223197e-10 lua=-2.906534191e-16 ub=1.485697036e-18 lub=3.071782747e-26 uc=2.621592345e-11 luc=-3.315325625e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.484334062e+00 la0=-1.032456821e-6 ags=3.532558268e-01 lags=-5.248898949e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.269093046e-02 lketa=8.872369085e-08 wketa=-1.734723476e-24 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=-3.606890755e-01 lpclm=3.532385178e-06 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=2.958440708e-03 lpdiblc2=1.526220364e-9 pdiblcb=-4.385714527e+00 lpdiblcb=1.723302489e-5 drout=0.56 pscbe1=7.776031919e+08 lpscbe1=-1.279409298e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912647966e-01 lkt1=-9.663152887e-9 kt2=-2.057567252e-02 lkt2=-4.849174381e-10 at=140000.0 ute=-1.487467585e+00 lute=1.588528060e-6 ua1=1.252925832e-09 lua1=8.005490075e-16 ub1=-9.359247047e-19 lub1=-4.878713775e-26 uc1=-3.045817068e-11 luc1=4.810766883e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.57 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.089124405e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.563726162e-8 k1=4.422672016e-01 lk1=1.896350346e-7 k2=1.499972931e-02 lk2=-9.125365600e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.664948260e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.651125123e-8 nfactor=3.266684827e+00 lnfactor=-1.647874417e-6 eta0=0.08 etab=-0.07 u0=2.967601883e-02 lu0=-3.669514476e-9 ua=-2.520500308e-10 lua=-1.769732966e-15 ub=9.297082108e-19 lub=2.227919503e-24 uc=-2.649083338e-12 luc=1.107557462e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.366787166e+00 la0=-5.679254763e-7 ags=2.093761749e-01 lags=5.161062732e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.791565865e-02 lketa=-7.174871712e-08 wketa=1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.098057438e-01 lpclm=9.229324121e-8 pdiblc1=0.39 pdiblc2=1.439337851e-03 lpdiblc2=7.529534081e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.917747749e+08 lpscbe1=2.112427606e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.956911592e-01 lkt1=7.829305460e-9 kt2=-2.362580522e-02 lkt2=1.156884401e-8 at=1.681070864e+05 lat=-1.110758607e-1 ute=-1.732577830e+00 lute=2.557174581e-6 ua1=-6.478469656e-10 lua1=8.312176910e-15 ub1=7.966432982e-19 lub1=-6.895689710e-24 pub1=-3.081487911e-45 uc1=-6.637324182e-12 luc1=-4.602948185e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.58 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.220559925e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.998261211e-8 k1=5.966824121e-01 lk1=-1.117650811e-7 k2=-4.993686404e-02 lk2=3.549484675e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.015830594e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.736268633e-8 nfactor=2.840858871e+00 lnfactor=-8.167128236e-7 eta0=1.537409836e-01 leta0=-1.439336249e-7 etab=-5.631671062e-02 letab=-2.670815255e-8 u0=2.951753534e-02 lu0=-3.360173574e-9 ua=-9.343234264e-10 lua=-4.380164887e-16 ub=1.955048112e-18 lub=2.265780315e-25 uc=3.881630995e-11 luc=2.982023293e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.048119000e+04 lvsat=1.857958438e-2 a0=1.413345773e+00 la0=-6.588023348e-7 ags=3.053090149e-01 lags=3.288567856e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.634123739e-02 lketa=3.415428738e-8 dwg=0.0 dwb=0.0 pclm=4.321841752e-01 lpclm=2.438013063e-7 pdiblc1=4.388270976e-01 lpdiblc1=-9.530468411e-8 pdiblc2=4.811682871e-03 lpdiblc2=9.471179099e-10 pdiblcb=-1.800242252e-03 lpdiblcb=-4.528316635e-8 drout=7.148712196e-01 ldrout=-3.022901909e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.114225720e-08 lalpha0=-2.229550126e-15 alpha1=9.956377930e-01 lalpha1=-2.842676410e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.250339102e-01 lkt1=6.510286367e-8 kt2=-6.229275676e-05 lkt2=-3.442432826e-8 at=1.354586873e+05 lat=-4.735007080e-2 ute=1.718178647e-01 lute=-1.159979192e-06 pute=4.440892099e-28 ua1=5.861327436e-09 lua1=-4.392956931e-15 ub1=-4.609958711e-18 lub1=3.657354026e-24 uc1=-7.616316627e-11 luc1=8.967668832e-17 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.59 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.788791820e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.106302280e-9 k1=4.031517729e-01 lk1=7.245305732e-8 k2=7.261457465e-03 lk2=-1.895114872e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.117788567e-01 ldsub=4.590079015e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.566723314e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.075744911e-9 nfactor=8.992262257e-01 lnfactor=1.031490401e-6 eta0=-4.380243872e-01 leta0=4.193565881e-07 weta0=9.714451465e-23 peta0=-8.673617380e-30 etab=-1.603474931e-01 letab=7.231677273e-8 u0=2.913828546e-02 lu0=-2.999172815e-9 ua=-1.313229939e-09 lua=-7.734257874e-17 ub=2.320380300e-18 lub=-1.211747371e-25 uc=6.345977625e-11 luc=6.362585589e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.815607246e+04 lvsat=2.079281959e-2 a0=1.742630488e-02 la0=6.699468839e-7 ags=2.491491296e-01 lags=3.823143134e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.675999412e-02 lketa=-3.542938598e-08 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=8.584974222e-01 lpclm=-1.619981737e-07 wpclm=-8.881784197e-22 pdiblc1=5.163711879e-01 lpdiblc1=-1.691174303e-07 wpdiblc1=4.440892099e-22 pdiblc2=9.603259256e-03 lpdiblc2=-3.613892611e-09 ppdiblc2=3.469446952e-30 pdiblcb=-7.139951550e-02 lpdiblcb=2.096705946e-8 drout=-1.473977191e-01 ldrout=5.184872287e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.771548560e-08 lalpha0=1.032328652e-15 alpha1=5.587244140e-01 lalpha1=1.316219031e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.438766302e-01 lkt1=-1.214920922e-8 kt2=-3.611529325e-02 lkt2=-1.061620977e-10 at=1.178750201e+05 lat=-3.061251210e-2 ute=-8.848952854e-01 lute=-1.541140217e-7 ua1=1.384291714e-09 lua1=-1.313516911e-16 ub1=-8.472332519e-19 lub1=7.568715372e-26 uc1=-1.072283955e-12 luc1=1.819910418e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.60 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.218604304e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.352871179e-8 k1=2.860351215e-01 lk1=1.253758469e-7 k2=4.425283035e-02 lk2=-3.566684729e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.960437946e-01 ldsub=5.301116574e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590352e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.187591359e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.205650776e-8 nfactor=3.662754514e+00 lnfactor=-2.172955256e-7 eta0=8.851262253e-01 leta0=-1.785500338e-7 etab=3.496458970e-02 letab=-1.594104657e-08 wetab=9.107298249e-24 petab=2.385244779e-30 u0=1.731479636e-02 lu0=2.343637264e-9 ua=-1.735371739e-09 lua=1.134152799e-16 ub=1.962422486e-18 lub=4.057959792e-26 uc=6.541098952e-11 luc=5.480869385e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.809020490e+04 lvsat=1.178496389e-2 a0=1.5 ags=9.701952848e-01 lags=5.648725571e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=9.946273253e-03 lketa=-1.879396498e-8 dwg=0.0 dwb=0.0 pclm=7.111109993e-01 lpclm=-9.539704948e-8 pdiblc1=-3.137998472e-02 lpdiblc1=7.840091731e-8 pdiblc2=-3.885586127e-03 lpdiblc2=2.481460330e-09 wpdiblc2=1.734723476e-24 ppdiblc2=4.336808690e-31 pdiblcb=3.822571337e-02 lpdiblcb=-2.857049858e-8 drout=1.401075642e+00 ldrout=-1.812384623e-7 pscbe1=8.069286528e+08 lpscbe1=-3.130926566e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.678320160e-08 lalpha0=-3.065199922e-15 alpha1=0.85 beta0=1.348853896e+01 lbeta0=1.678561862e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.948281184e-01 lkt1=1.087480021e-8 kt2=-4.238347137e-02 lkt2=2.726308500e-9 at=6.741939690e+04 lat=-7.812574629e-3 ute=-1.150766511e+00 lute=-3.397186617e-8 ua1=1.995991029e-09 lua1=-4.077669889e-16 ub1=-1.800173492e-18 lub1=5.063027425e-25 wub1=7.703719778e-40 uc1=-4.799819162e-11 luc1=3.940403026e-17 puc1=-1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.61 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='1.095288763e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.191048969e-07 wvth0=-4.787991876e-07 pvth0=9.666045880e-14 k1=0.90707349 k2=-3.926179182e-01 lk2=5.252905629e-08 wk2=2.232236364e-07 pk2=-4.506461094e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586393070e-01 ldsub=-1.878912639e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.237493850e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907129e-8 nfactor=-5.074445767e+00 lnfactor=1.546579204e-06 wnfactor=9.063478171e-06 pnfactor=-1.829744037e-12 eta0=6.941422985e-04 leta0=-4.640229594e-16 etab=-0.043998 u0=5.426925210e-02 lu0=-5.116765215e-09 wu0=-2.108319836e-08 pu0=4.256297168e-15 ua=-1.410310372e-09 lua=4.779156618e-17 wua=2.086995943e-16 pua=-4.213248280e-23 ub=3.629264811e-18 lub=-2.959241974e-25 wub=-1.461354754e-24 pub=2.950197592e-31 uc=3.259345894e-10 luc=-4.711389547e-17 wuc=-2.669421929e-16 puc=5.389055684e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.042030007e+05 lvsat=-1.165600343e-02 wvsat=-7.414857538e-02 pvsat=1.496918855e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.227757627e-01 lketa=8.875249237e-08 wketa=3.569235300e-07 pketa=-7.205607915e-14 dwg=0.0 dwb=0.0 pclm=3.406610229e-01 lpclm=-2.061023780e-08 wpclm=1.032332671e-07 ppclm=-2.084083520e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.517434155e-08 lalpha0=1.549928085e-14 walpha0=7.687583723e-14 palpha0=-1.551977089e-20 alpha1=0.85 beta0=1.687431802e+01 lbeta0=-5.156682759e-07 wbeta0=-2.104933638e-06 pbeta0=4.249461078e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.237567913e-01 lkt1=3.690304963e-08 wkt1=1.830377077e-07 pkt1=-3.695183546e-14 kt2=-0.028878939 at=1.512280812e+05 lat=-2.473195562e-02 wat=-1.830377077e-01 pat=3.695183546e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.62 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-5.105009820e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.266826037e-08 wvth0=1.140425525e-06 pvth0=-1.168845155e-13 k1=0.90707349 k2=2.973095529e-01 lk2=-3.845926853e-08 wk2=-4.863109625e-07 pk2=4.850952149e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.595374184e+01 lnfactor=-2.545449205e-06 wnfactor=-2.915563694e-05 pnfactor=3.210631083e-12 eta0=0.00069413878 etab=-0.043998 u0=-1.562949565e-02 lu0=4.101551537e-09 wu0=5.041818816e-08 pu0=-5.173377188e-15 ua=-7.661145631e-10 lua=-3.716562134e-17 wua=-4.662293085e-16 pua=4.687781583e-23 ub=-1.679499335e-18 lub=4.042009269e-25 wub=4.641474923e-24 pub=-5.098275216e-31 uc=-4.127972759e-10 luc=5.031080165e-17 wuc=6.228651167e-16 puc=-6.345812096e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.771363641e+04 lvsat=3.706730415e-03 wvsat=7.480820510e-02 pvsat=-4.675380620e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.602767334e-01 lketa=-6.726965388e-08 wketa=-8.328215699e-07 pketa=8.484869437e-14 dwg=0.0 dwb=0.0 pclm=1.843819698e-01 wpclm=-5.479431229e-8 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.722134503e-07 lalpha0=-1.448884853e-14 walpha0=-1.793769535e-13 palpha0=1.827510340e-20 alpha1=0.85 beta0=9.956060290e+00 lbeta0=3.967184716e-07 wbeta0=4.911511823e-06 pbeta0=-5.003897360e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=1.176427130e-01 lkt1=-3.449725840e-08 wkt1=-4.270879846e-07 pkt1=4.351215096e-14 kt2=-0.028878939 at=-2.978829660e+05 lat=3.449725840e-02 wat=4.270879846e-01 pat=-4.351215096e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.63 nmos lmin=2.0e-05 lmax=0.0001 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.381335181e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.405355939e-06 wvth0=4.549834204e-08 pvth0=-4.547644869e-12 k1=7.154905561e-01 lk1=-1.474118689e-05 wk1=-1.240805547e-07 pk1=1.240208483e-11 k2=-1.016607536e-01 lk2=6.193539053e-06 wk2=5.213269236e-08 pk2=-5.210760663e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.033776573e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.897824770e-07 wvoff=-4.122631500e-09 pvoff=4.120647731e-13 nfactor=3.186706537e+00 lnfactor=-3.039602036e-05 wnfactor=-2.558515196e-07 pnfactor=2.557284064e-11 eta0=0.08 etab=-0.07 u0=2.200495044e-02 lu0=4.644113787e-07 wu0=3.909076108e-09 pu0=-3.907195099e-13 ua=-1.673038924e-09 lua=6.153965584e-14 wua=5.179959178e-16 pua=-5.177466633e-20 ub=2.292094659e-18 lub=-4.889072887e-23 wub=-4.115264804e-25 pub=4.113284580e-29 uc=8.402650129e-11 luc=-3.547242409e-15 wuc=-2.985809820e-17 puc=2.984373078e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.375248734e+00 la0=-1.264264776e-06 wa0=-1.064165836e-08 pa0=1.063653770e-12 ags=3.421095776e-01 lags=2.769089311e-07 wags=2.330817324e-09 pags=-2.329695758e-13 a1=0.0 a2=0.42385546 b0=1.625315014e-07 lb0=-9.901483353e-12 wb0=-8.334346181e-14 pb0=8.330335777e-18 b1=6.451682942e-09 lb1=-3.930390767e-13 wb1=-3.308316149e-15 pb1=3.306724221e-19 keta=-9.249672675e-03 lketa=4.700809603e-07 wketa=3.956798509e-09 pketa=-3.954894537e-13 dwg=0.0 dwb=0.0 pclm=-8.716177534e-02 lpclm=1.039867139e-05 wpclm=8.752842790e-08 ppclm=-8.748631010e-12 pdiblc1=0.39 pdiblc2=-2.457898125e-03 lpdiblc2=3.416580769e-07 wpdiblc2=2.875828386e-09 ppdiblc2=-2.874444566e-13 pdiblcb=3.398697693e+00 lpdiblcb=-3.422050243e-04 wpdiblcb=-2.880432190e-06 ppdiblcb=2.879046155e-10 drout=0.56 pscbe1=-6.123914678e+08 lpscbe1=8.369885234e+04 wpscbe1=7.045158645e+02 ppscbe1=-7.041768585e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.768591117e-01 lkt1=-9.516306930e-07 wkt1=-8.010132774e-09 pkt1=8.006278379e-13 kt2=-4.337984021e-02 lkt2=1.385523899e-06 wkt2=1.166232918e-08 pkt2=-1.165671738e-12 at=2.296280475e+05 lat=-5.460176107e+00 wat=-4.595977821e-02 pat=4.593766283e-6 ute=-8.464739260e-01 lute=-2.687966695e-05 wute=-2.262534225e-07 pute=2.261445516e-11 ua1=7.579576041e-10 lua1=3.628677036e-14 wua1=3.054355546e-16 pua1=-3.052885821e-20 ub1=1.206897810e-20 lub1=-5.812591474e-23 wub1=-4.892615361e-25 pub1=4.890261084e-29 uc1=1.246986510e-10 luc1=-9.083655835e-15 wuc1=-7.645958654e-17 puc1=7.642279495e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.64 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='8.297835176e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.408798246e-06 wvth0=-3.033222803e-07 pvth0=2.411982677e-12 k1=-3.525955983e-01 lk1=6.569140963e-06 wk1=8.272036978e-07 pk1=-6.577825368e-12 k2=3.470977731e-01 lk2=-2.760037669e-06 wk2=-3.475512824e-07 pk2=2.763686439e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.388652938e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.182626241e-07 wvoff=2.748421000e-08 pvoff=-2.185511673e-13 nfactor=9.843351301e-01 lnfactor=1.354543186e-05 wnfactor=1.705676798e-06 pnfactor=-1.356333892e-11 eta0=0.08 etab=-0.07 u0=5.565430088e-02 lu0=-2.069564571e-07 wu0=-2.606050738e-08 pu0=2.072300535e-13 ua=2.785873025e-09 lua=-2.742402475e-14 wua=-3.453306118e-15 pua=2.746027931e-20 ub=-1.250327738e-18 lub=2.178726124e-23 wub=2.743509869e-24 pub=-2.181606400e-29 uc=-1.729921861e-10 luc=1.580763855e-15 wuc=1.990539880e-16 puc=-1.582853625e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.283645276e+00 la0=5.633965293e-07 wa0=7.094438908e-08 pa0=-5.641413395e-13 ags=3.621732670e-01 lags=-1.233994126e-07 wags=-1.553878216e-08 pags=1.235625466e-13 a1=0.0 a2=0.42385546 b0=-5.548895148e-07 lb0=4.412415390e-12 wb0=5.556230788e-13 pb0=-4.418248603e-18 b1=-2.202632220e-08 lb1=1.751506930e-13 wb1=2.205544100e-14 pb1=-1.753822422e-19 keta=2.481047248e-02 lketa=-2.094830027e-07 wketa=-2.637865673e-08 pketa=2.097599392e-13 dwg=0.0 dwb=0.0 pclm=6.662834539e-01 lpclm=-4.633978166e-06 wpclm=-5.835228527e-07 ppclm=4.640104285e-12 pdiblc1=0.39 pdiblc2=2.229724977e-02 lpdiblc2=-1.522536880e-07 wpdiblc2=-1.917218924e-08 ppdiblc2=1.524549673e-13 pdiblcb=-2.139607977e+01 lpdiblcb=1.524974251e-04 wpdiblcb=1.920288127e-05 ppdiblcb=-1.526990267e-10 drout=0.56 pscbe1=5.452085294e+09 lpscbe1=-3.729886634e+04 wpscbe1=-4.696772430e+03 ppscbe1=3.734817545e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.458103824e-01 lkt1=4.240768545e-07 wkt1=5.340088516e-08 pkt1=-4.246374841e-13 kt2=5.700955888e-02 lkt2=-6.174334449e-07 wkt2=-7.774886118e-08 pkt2=6.182496920e-13 at=-1.659939974e+05 lat=2.433227854e+00 wat=3.063985214e-01 pat=-2.436444581e-6 ute=-2.794064736e+00 lute=1.197843312e-05 wute=1.508356150e-06 pute=-1.199426861e-11 ua1=3.387148680e-09 lua1=-1.617053711e-14 wua1=-2.036237031e-15 pua1=1.619191456e-20 ub1=-4.199497242e-18 lub1=2.590275331e-23 wub1=3.261743574e-24 pub1=-2.593699675e-29 uc1=-5.334659258e-10 luc1=4.047965479e-15 wuc1=5.097305769e-16 puc1=-4.053316890e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.65 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.256857190e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.351260879e-9 k1=4.569800848e-01 lk1=1.314914708e-7 k2=8.004757165e-03 lk2=-6.361035850e-08 wk2=2.175180609e-24 pk2=-1.764539036e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.167594931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.247992715e-8 nfactor=2.527768098e+00 lnfactor=1.272236568e-6 eta0=0.08 etab=-0.07 u0=3.049833504e-02 lu0=-6.919210278e-9 ua=-6.263223197e-10 lua=-2.906534191e-16 ub=1.485697036e-18 lub=3.071782747e-26 uc=2.621592345e-11 luc=-3.315325625e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.484334062e+00 la0=-1.032456821e-6 ags=3.532558268e-01 lags=-5.248898949e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.269093046e-02 lketa=8.872369085e-08 wketa=-6.938893904e-24 dwg=0.0 dwb=0.0 pclm=-3.606890755e-01 lpclm=3.532385178e-06 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=2.958440708e-03 lpdiblc2=1.526220364e-9 pdiblcb=-4.385714527e+00 lpdiblcb=1.723302489e-5 drout=0.56 pscbe1=7.776031919e+08 lpscbe1=-1.279409298e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912647966e-01 lkt1=-9.663152887e-9 kt2=-2.057567252e-02 lkt2=-4.849174381e-10 at=140000.0 ute=-1.487467585e+00 lute=1.588528060e-6 ua1=1.252925832e-09 lua1=8.005490075e-16 ub1=-9.359247047e-19 lub1=-4.878713775e-26 uc1=-3.045817068e-11 luc1=4.810766883e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.66 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.089124405e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.563726162e-8 k1=4.422672016e-01 lk1=1.896350346e-7 k2=1.499972931e-02 lk2=-9.125365600e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.664948260e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.651125123e-8 nfactor=3.266684827e+00 lnfactor=-1.647874417e-06 wnfactor=-3.552713679e-21 eta0=0.08 etab=-0.07 u0=2.967601883e-02 lu0=-3.669514476e-9 ua=-2.520500308e-10 lua=-1.769732966e-15 ub=9.297082108e-19 lub=2.227919503e-24 uc=-2.649083338e-12 luc=1.107557462e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.366787166e+00 la0=-5.679254763e-7 ags=2.093761749e-01 lags=5.161062732e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.791565865e-02 lketa=-7.174871712e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.098057438e-01 lpclm=9.229324121e-8 pdiblc1=0.39 pdiblc2=1.439337851e-03 lpdiblc2=7.529534081e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.917747749e+08 lpscbe1=2.112427606e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.956911592e-01 lkt1=7.829305460e-9 kt2=-2.362580522e-02 lkt2=1.156884401e-8 at=1.681070864e+05 lat=-1.110758607e-1 ute=-1.732577830e+00 lute=2.557174581e-6 ua1=-6.478469656e-10 lua1=8.312176910e-15 pua1=3.308722450e-36 ub1=7.966432982e-19 lub1=-6.895689710e-24 uc1=-6.637324182e-12 luc1=-4.602948185e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.67 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.220559925e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.998261211e-8 k1=5.966824121e-01 lk1=-1.117650811e-7 k2=-4.993686404e-02 lk2=3.549484675e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-07 wdsub=8.881784197e-22 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.015830594e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.736268633e-8 nfactor=2.840858871e+00 lnfactor=-8.167128236e-7 eta0=1.537409836e-01 leta0=-1.439336249e-7 etab=-5.631671062e-02 letab=-2.670815255e-8 u0=2.951753534e-02 lu0=-3.360173574e-9 ua=-9.343234264e-10 lua=-4.380164887e-16 ub=1.955048112e-18 lub=2.265780315e-25 uc=3.881630995e-11 luc=2.982023293e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.048119000e+04 lvsat=1.857958438e-2 a0=1.413345773e+00 la0=-6.588023348e-7 ags=3.053090149e-01 lags=3.288567856e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.634123739e-02 lketa=3.415428738e-08 wketa=1.387778781e-23 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=4.321841752e-01 lpclm=2.438013063e-7 pdiblc1=4.388270976e-01 lpdiblc1=-9.530468411e-8 pdiblc2=4.811682871e-03 lpdiblc2=9.471179099e-10 pdiblcb=-1.800242252e-03 lpdiblcb=-4.528316635e-8 drout=7.148712196e-01 ldrout=-3.022901909e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.114225720e-08 lalpha0=-2.229550126e-15 alpha1=9.956377930e-01 lalpha1=-2.842676410e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.250339102e-01 lkt1=6.510286367e-8 kt2=-6.229275676e-05 lkt2=-3.442432826e-8 at=1.354586873e+05 lat=-4.735007080e-2 ute=1.718178647e-01 lute=-1.159979192e-6 ua1=5.861327436e-09 lua1=-4.392956931e-15 ub1=-4.609958711e-18 lub1=3.657354026e-24 pub1=-3.081487911e-45 uc1=-7.616316627e-11 luc1=8.967668832e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.68 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.788791820e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.106302280e-9 k1=4.031517729e-01 lk1=7.245305732e-8 k2=7.261457465e-03 lk2=-1.895114872e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.117788567e-01 ldsub=4.590079015e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.566723314e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.075744911e-9 nfactor=8.992262257e-01 lnfactor=1.031490401e-6 eta0=-4.380243872e-01 leta0=4.193565881e-07 weta0=2.081668171e-22 peta0=-1.561251128e-28 etab=-1.603474931e-01 letab=7.231677273e-8 u0=2.913828546e-02 lu0=-2.999172815e-9 ua=-1.313229939e-09 lua=-7.734257874e-17 ub=2.320380300e-18 lub=-1.211747371e-25 uc=6.345977625e-11 luc=6.362585589e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.815607246e+04 lvsat=2.079281959e-2 a0=1.742630488e-02 la0=6.699468839e-7 ags=2.491491296e-01 lags=3.823143134e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.675999412e-02 lketa=-3.542938598e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=8.584974222e-01 lpclm=-1.619981737e-7 pdiblc1=5.163711879e-01 lpdiblc1=-1.691174303e-7 pdiblc2=9.603259256e-03 lpdiblc2=-3.613892611e-9 pdiblcb=-7.139951550e-02 lpdiblcb=2.096705946e-08 wpdiblcb=5.551115123e-23 drout=-1.473977191e-01 ldrout=5.184872287e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.771548560e-08 lalpha0=1.032328652e-15 alpha1=5.587244140e-01 lalpha1=1.316219031e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.438766302e-01 lkt1=-1.214920922e-8 kt2=-3.611529325e-02 lkt2=-1.061620977e-10 at=1.178750201e+05 lat=-3.061251210e-2 ute=-8.848952854e-01 lute=-1.541140217e-7 ua1=1.384291714e-09 lua1=-1.313516911e-16 ub1=-8.472332519e-19 lub1=7.568715372e-26 uc1=-1.072283955e-12 luc1=1.819910418e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.69 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.218604304e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.352871179e-8 k1=2.860351215e-01 lk1=1.253758469e-7 k2=4.425283035e-02 lk2=-3.566684729e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.960437946e-01 ldsub=5.301116574e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590352e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.187591359e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.205650776e-8 nfactor=3.662754514e+00 lnfactor=-2.172955256e-07 wnfactor=-3.552713679e-21 eta0=8.851262253e-01 leta0=-1.785500338e-7 etab=3.496458970e-02 letab=-1.594104657e-08 wetab=-7.806255642e-24 petab=1.192622390e-30 u0=1.731479636e-02 lu0=2.343637264e-9 ua=-1.735371739e-09 lua=1.134152799e-16 ub=1.962422486e-18 lub=4.057959792e-26 uc=6.541098952e-11 luc=5.480869385e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.809020490e+04 lvsat=1.178496389e-2 a0=1.5 ags=9.701952848e-01 lags=5.648725571e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=9.946273253e-03 lketa=-1.879396498e-08 pketa=6.938893904e-30 dwg=0.0 dwb=0.0 pclm=7.111109993e-01 lpclm=-9.539704948e-8 pdiblc1=-3.137998472e-02 lpdiblc1=7.840091731e-8 pdiblc2=-3.885586127e-03 lpdiblc2=2.481460330e-09 wpdiblc2=1.734723476e-24 ppdiblc2=-8.673617380e-31 pdiblcb=3.822571337e-02 lpdiblcb=-2.857049858e-08 ppdiblcb=6.938893904e-30 drout=1.401075642e+00 ldrout=-1.812384623e-7 pscbe1=8.069286528e+08 lpscbe1=-3.130926566e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.678320160e-08 lalpha0=-3.065199922e-15 alpha1=0.85 beta0=1.348853896e+01 lbeta0=1.678561862e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.948281184e-01 lkt1=1.087480021e-8 kt2=-4.238347137e-02 lkt2=2.726308500e-9 at=6.741939690e+04 lat=-7.812574629e-3 ute=-1.150766511e+00 lute=-3.397186617e-8 ua1=1.995991029e-09 lua1=-4.077669889e-16 ub1=-1.800173492e-18 lub1=5.063027425e-25 wub1=-7.703719778e-40 uc1=-4.799819162e-11 luc1=3.940403026e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.70 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.171217118e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.257205455e-8 k1=0.90707349 k2=-1.696889938e-01 lk2=7.523942113e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586393070e-01 ldsub=-1.878912639e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.237493850e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907129e-8 nfactor=3.977066305e+00 lnfactor=-2.807491043e-7 eta0=6.941422985e-04 leta0=-4.640229594e-16 etab=-0.043998 u0=3.321388893e-02 lu0=-8.660874433e-10 ua=-1.201886315e-09 lua=5.714708987e-18 ub=2.169839417e-18 lub=-1.293939433e-27 uc=5.934482814e-11 luc=6.705512110e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.301523203e+05 lvsat=3.293421972e-3 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.663234627e-01 lketa=1.679154558e-8 dwg=0.0 dwb=0.0 pclm=4.437579959e-01 lpclm=-4.142355779e-8 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.16e-8 alpha1=0.85 beta0=1.477216343e+01 lbeta0=-9.128320512e-8 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.24096074 kt2=-0.028878939 at=-3.156797014e+04 lat=1.217109402e-2 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.71 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='3.387388291e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.414135840e-08 wvth0=2.900630188e-07 pvth0=-3.825380098e-14 k1=0.90707349 k2=-2.073415957e-01 lk2=1.248960491e-08 wk2=1.900733504e-08 pk2=-2.506706352e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587132747e-01 ldsub=-1.163384807e-11 wdsub=-8.833135943e-11 pdsub=1.164922801e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-1.647025640e+01 lnfactor=2.415864262e-06 wnfactor=1.332444583e-05 pnfactor=-1.757241241e-12 eta0=-1.170125918e-02 leta0=1.634717632e-09 weta0=1.241178584e-08 peta0=-1.636878729e-15 etab=-0.043998 u0=2.921138503e-02 lu0=-3.382332261e-10 wu0=5.518027838e-09 pu0=-7.277230293e-16 ua=-2.224465580e-09 lua=1.405734851e-16 wua=9.940496487e-16 pua=-1.310962617e-22 ub=6.672116778e-18 lub=-5.950587801e-25 wub=-3.721182026e-24 pub=4.907532068e-31 uc=1.374951311e-10 luc=-3.601028000e-18 wuc=7.184522311e-17 puc=-9.475019870e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.027263399e+05 lvsat=6.910387687e-03 wvsat=5.977565477e-02 pvsat=-7.883273127e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.535906376e-01 lketa=8.105282788e-08 wketa=4.827827337e-07 pketa=-6.366986971e-14 dwg=0.0 dwb=0.0 pclm=1.014455691e-01 lpclm=3.720947357e-09 wpclm=2.825173034e-08 ppclm=-3.725866449e-15 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.926680000e-09 lalpha0=3.762127085e-15 alpha1=0.85 beta0=1.843253461e+01 lbeta0=-5.740166171e-07 wbeta0=-3.576168398e-06 pbeta0=4.716286645e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-6.660261012e-01 lkt1=5.605804490e-08 wkt1=3.576168398e-07 pkt1=-4.716286645e-14 kt2=-0.028878939 at=3.607852051e+05 lat=-3.957283509e-02 wat=-2.324509459e-01 pat=3.065586319e-8 ute=-4.261814637e-01 lute=-1.177514986e-07 wute=-8.940420995e-07 pute=1.179071661e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.72 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.73 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.692529713e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.580977549e-7 k1=6.306233093e-01 lk1=-1.249298787e-6 k2=-6.600361066e-02 lk2=5.248953755e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.061974093e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.150850668e-8 nfactor=3.011712041e+00 lnfactor=-2.576028081e-6 eta0=0.08 etab=-0.07 u0=2.467863712e-02 lu0=3.935833502e-8 ua=-1.318745799e-09 lua=5.215415691e-15 ub=2.010623324e-18 lub=-4.143433547e-24 uc=6.360448918e-11 luc=-3.006247511e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.367970170e+00 la0=-1.071449988e-07 wa0=-1.776356839e-21 ags=3.437037843e-01 lags=2.346771630e-8 a1=0.0 a2=0.42385546 b0=1.055271613e-07 lb0=-8.391394287e-13 b1=4.188897416e-09 lb1=-3.330961377e-14 keta=-6.543345349e-03 lketa=3.983882560e-8 dwg=0.0 dwb=0.0 pclm=-2.729504833e-02 lpclm=8.812755480e-07 ppclm=2.220446049e-28 pdiblc1=0.39 pdiblc2=-4.909208011e-04 lpdiblc2=2.895513261e-8 pdiblcb=1.428571509e+00 lpdiblcb=-2.900148578e-05 wpdiblcb=1.110223025e-22 ppdiblcb=-3.108624469e-27 drout=0.56 pscbe1=-1.305244910e+08 lpscbe1=7.093382338e+03 ppscbe1=-3.814697266e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.823377938e-01 lkt1=-8.064961658e-8 kt2=-3.540316915e-02 lkt2=1.174215713e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.001224242e+00 lute=-2.278021137e-6 ua1=9.668660399e-10 lua1=3.075262429e-15 ub1=-3.225707215e-19 lub1=-4.926105023e-24 uc1=7.240266785e-11 luc1=-7.698294787e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.74 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.256857190e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.351260879e-9 k1=4.569800848e-01 lk1=1.314914708e-7 k2=8.004757165e-03 lk2=-6.361035850e-08 wk2=4.607859233e-25 pk2=9.486769009e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.167594931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.247992715e-8 nfactor=2.527768098e+00 lnfactor=1.272236568e-6 eta0=0.08 etab=-0.07 u0=3.049833504e-02 lu0=-6.919210278e-9 ua=-6.263223197e-10 lua=-2.906534191e-16 ub=1.485697036e-18 lub=3.071782747e-26 uc=2.621592345e-11 luc=-3.315325625e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.484334062e+00 la0=-1.032456821e-6 ags=3.532558268e-01 lags=-5.248898949e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.269093046e-02 lketa=8.872369085e-08 wketa=6.938893904e-24 pketa=-4.163336342e-29 dwg=0.0 dwb=0.0 pclm=-3.606890755e-01 lpclm=3.532385178e-06 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=2.958440708e-03 lpdiblc2=1.526220364e-9 pdiblcb=-4.385714527e+00 lpdiblcb=1.723302489e-5 drout=0.56 pscbe1=7.776031919e+08 lpscbe1=-1.279409298e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912647966e-01 lkt1=-9.663152887e-9 kt2=-2.057567252e-02 lkt2=-4.849174381e-10 at=140000.0 ute=-1.487467585e+00 lute=1.588528060e-6 ua1=1.252925832e-09 lua1=8.005490075e-16 ub1=-9.359247047e-19 lub1=-4.878713775e-26 uc1=-3.045817068e-11 luc1=4.810766883e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.75 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.089124405e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.563726162e-8 k1=4.422672016e-01 lk1=1.896350346e-7 k2=1.499972931e-02 lk2=-9.125365600e-08 pk2=2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.664948260e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.651125123e-8 nfactor=3.266684827e+00 lnfactor=-1.647874417e-6 eta0=0.08 etab=-0.07 u0=2.967601883e-02 lu0=-3.669514476e-9 ua=-2.520500308e-10 lua=-1.769732966e-15 ub=9.297082108e-19 lub=2.227919503e-24 uc=-2.649083338e-12 luc=1.107557462e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.366787166e+00 la0=-5.679254763e-07 wa0=-1.776356839e-21 ags=2.093761749e-01 lags=5.161062732e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.791565865e-02 lketa=-7.174871712e-8 dwg=0.0 dwb=0.0 pclm=5.098057438e-01 lpclm=9.229324121e-8 pdiblc1=0.39 pdiblc2=1.439337851e-03 lpdiblc2=7.529534081e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.917747749e+08 lpscbe1=2.112427606e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.956911592e-01 lkt1=7.829305460e-9 kt2=-2.362580522e-02 lkt2=1.156884401e-8 at=1.681070864e+05 lat=-1.110758607e-1 ute=-1.732577830e+00 lute=2.557174581e-6 ua1=-6.478469656e-10 lua1=8.312176910e-15 ub1=7.966432982e-19 lub1=-6.895689710e-24 uc1=-6.637324182e-12 luc1=-4.602948185e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.76 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.220559925e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.998261211e-8 k1=5.966824121e-01 lk1=-1.117650811e-7 k2=-4.993686404e-02 lk2=3.549484675e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.015830594e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.736268633e-8 nfactor=2.840858871e+00 lnfactor=-8.167128236e-7 eta0=1.537409836e-01 leta0=-1.439336249e-7 etab=-5.631671062e-02 letab=-2.670815255e-8 u0=2.951753534e-02 lu0=-3.360173574e-9 ua=-9.343234264e-10 lua=-4.380164887e-16 ub=1.955048112e-18 lub=2.265780315e-25 uc=3.881630995e-11 luc=2.982023293e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.048119000e+04 lvsat=1.857958438e-2 a0=1.413345773e+00 la0=-6.588023348e-7 ags=3.053090149e-01 lags=3.288567856e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.634123739e-02 lketa=3.415428738e-8 dwg=0.0 dwb=0.0 pclm=4.321841752e-01 lpclm=2.438013063e-7 pdiblc1=4.388270976e-01 lpdiblc1=-9.530468411e-8 pdiblc2=4.811682871e-03 lpdiblc2=9.471179099e-10 pdiblcb=-1.800242252e-03 lpdiblcb=-4.528316635e-8 drout=7.148712196e-01 ldrout=-3.022901909e-07 wdrout=-8.881784197e-22 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.114225720e-08 lalpha0=-2.229550126e-15 alpha1=9.956377930e-01 lalpha1=-2.842676410e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.250339102e-01 lkt1=6.510286367e-8 kt2=-6.229275676e-05 lkt2=-3.442432826e-8 at=1.354586873e+05 lat=-4.735007080e-2 ute=1.718178647e-01 lute=-1.159979192e-6 ua1=5.861327436e-09 lua1=-4.392956931e-15 ub1=-4.609958711e-18 lub1=3.657354026e-24 uc1=-7.616316627e-11 luc1=8.967668832e-17 wuc1=-5.169878828e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.77 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='3.776701875e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.874207165e-07 wvth0=1.692815536e-07 pvth0=-1.611358945e-13 k1=-1.898082116e-01 lk1=6.368804003e-07 wk1=4.988702801e-07 pk1=-4.748651411e-13 k2=1.537496906e-01 lk2=-1.583905145e-07 wk2=-1.232437733e-07 pk2=1.173134061e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.913519444e-01 ldsub=6.534477978e-08 wdsub=1.718561065e-08 pdsub=-1.635865625e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.445898026e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.425384674e-09 wvoff=-1.016529729e-08 pvoff=9.676153345e-15 nfactor=-7.611517243e-01 lnfactor=2.611972624e-06 wnfactor=1.396912498e-06 pnfactor=-1.329694465e-12 eta0=-4.380243871e-01 leta0=4.193565880e-07 weta0=-1.131280035e-16 peta0=1.076843614e-22 etab=-1.624411764e-01 letab=7.430971005e-08 wetab=1.761461792e-09 petab=-1.676702012e-15 u0=4.593331033e-02 lu0=-1.898603789e-08 wu0=-1.413002392e-08 pu0=1.345010129e-14 ua=-1.068396291e-09 lua=-3.103950768e-16 wua=-2.059839347e-16 pua=1.960721937e-22 ub=2.641676602e-18 lub=-4.270105826e-25 wub=-2.703136476e-25 pub=2.573064252e-31 uc=-1.040549865e-10 luc=1.658167055e-16 wuc=1.409338552e-16 puc=-1.341522590e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.093215885e+05 lvsat=-2.087680530e-01 wvsat=-2.028978543e-01 pvsat=1.931346124e-7 a0=-7.557290596e-01 la0=1.405898785e-06 wa0=6.504726176e-07 pa0=-6.191725257e-13 ags=-6.041615430e+00 lags=6.370373573e-06 wags=5.292558621e-06 pags=-5.037885992e-12 a1=0.0 a2=0.42385546 b0=-3.959107428e-16 lb0=3.768599137e-22 wb0=3.330884179e-22 pb0=-3.170605363e-28 b1=1.061688972e-17 lb1=-1.010601560e-23 wb1=-8.932222891e-24 pb1=8.502413257e-30 keta=2.111120015e-01 lketa=-1.918729392e-07 wketa=-1.382729596e-07 pketa=1.316194030e-13 dwg=0.0 dwb=0.0 pclm=5.356347075e-01 lpclm=1.453287101e-07 wpclm=2.716315049e-07 ppclm=-2.585608685e-13 pdiblc1=-2.144901472e-01 lpdiblc1=5.265755882e-07 wpdiblc1=6.148897202e-07 ppdiblc1=-5.853018417e-13 pdiblc2=-8.442433845e-04 lpdiblc2=6.330886650e-09 wpdiblc2=8.789713817e-09 ppdiblc2=-8.366761578e-15 pdiblcb=-5.377395641e-01 lpdiblcb=4.648672912e-07 wpdiblcb=3.923421423e-07 ppdiblcb=-3.734630308e-13 drout=-1.473983893e-01 ldrout=5.184878667e-07 wdrout=5.638491238e-13 pdrout=-5.367172680e-19 pscbe1=-1.632377531e+09 lpscbe1=2.315333957e+03 wpscbe1=2.046412729e+03 ppscbe1=-1.947941395e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.595588937e-05 lalpha0=-2.467950376e-11 walpha0=-2.181394311e-11 palpha0=2.076427798e-17 alpha1=5.587244140e-01 lalpha1=1.316219031e-7 beta0=4.171771239e+01 lbeta0=-2.651722713e-05 wbeta0=-2.343730631e-05 pbeta0=2.230952656e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.987283855e-01 lkt1=4.006313448e-08 wkt1=4.614798848e-08 pkt1=-4.392739342e-14 kt2=-3.858331371e-02 lkt2=2.243099687e-09 wkt2=2.076399911e-09 pkt2=-1.976485623e-15 at=-1.465999106e+05 lat=2.211361494e-01 wat=2.225085777e-01 pat=-2.118016874e-7 ute=-1.449912404e+00 lute=3.837150378e-07 wute=4.753613319e-07 pute=-4.524874199e-13 ua1=-3.706807192e-10 lua1=1.539173224e-15 wua1=1.476496918e-15 pua1=-1.405449363e-21 ub1=-5.265767783e-19 lub1=-2.295396510e-25 wub1=-2.697753457e-25 pub1=2.567940258e-31 uc1=-2.252564936e-10 luc1=2.315957939e-16 wuc1=1.886111077e-16 puc1=-1.795353298e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.78 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='8.700280595e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.506645099e-08 wvth0=-2.087888861e-07 pvth0=9.706953816e-15 k1=1.471955090e+00 lk1=-1.140388620e-07 wk1=-9.977405595e-07 pk1=2.014248617e-13 k2=-2.631093814e-01 lk2=2.998017976e-08 wk2=2.585905907e-07 pk2=-5.523028809e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.368976191e-01 ldsub=4.476355475e-08 wdsub=-3.437122139e-08 pdsub=6.938896572e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590345e-03 lcdscd=-1.221701109e-09 wcdscd=6.181943846e-18 pcdscd=-2.793501541e-24 cit=0.0 voff='-1.429241933e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.178041876e-09 wvoff=2.033059438e-08 pvoff=-4.104360677e-15 nfactor=6.983510415e+00 lnfactor=-8.876930482e-07 wnfactor=-2.793824997e-06 pnfactor=5.640201845e-13 eta0=8.851262253e-01 leta0=-1.785500339e-07 weta0=-4.574474133e-17 peta0=7.723532924e-23 etab=3.915195620e-02 letab=-1.678639630e-08 wetab=-3.522923554e-09 petab=7.112113226e-16 u0=-8.847386534e-03 lu0=5.768318195e-09 wu0=2.201082003e-08 pu0=-2.881259410e-15 ua=-2.225039032e-09 lua=2.122698020e-16 wua=4.119678668e-16 pua=-8.316848429e-23 ub=1.319829883e-18 lub=1.703068349e-25 wub=5.406272940e-25 pub=-1.091423784e-31 uc=4.004405151e-10 luc=-6.215522629e-17 wuc=-2.818677105e-16 puc=5.690373529e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.659612950e+05 lvsat=9.637945173e-02 wvsat=3.820035160e-01 pvsat=-7.117120370e-8 a0=3.046310727e+00 la0=-3.121707552e-07 wa0=-1.300945233e-06 pa0=2.626361241e-13 ags=1.355172440e+01 lags=-2.483484424e-06 wags=-1.058511724e-05 pags=2.136934054e-12 a1=0.0 a2=0.42385546 b0=7.918214855e-16 lb0=-1.598537133e-22 wb0=-6.661768359e-22 pb0=1.344884458e-28 b1=-2.123377943e-17 lb1=4.286696626e-24 wb1=1.786444578e-23 pb1=-3.606492179e-30 keta=-3.187577415e-01 lketa=4.756513022e-08 wketa=2.765459191e-07 pketa=-5.582936669e-14 dwg=0.0 dwb=0.0 pclm=1.356836429e+00 lpclm=-2.257567451e-07 wpclm=-5.432630101e-07 ppclm=1.096744798e-13 pdiblc1=1.430342686e+00 lpdiblc1=-2.166931173e-07 wpdiblc1=-1.229779441e-06 ppdiblc1=2.482691034e-13 pdiblc2=1.700941914e-02 lpdiblc2=-1.736844226e-09 wpdiblc2=-1.757942762e-08 ppdiblc2=3.548952426e-15 pdiblcb=9.709058105e-01 lpdiblcb=-2.168608893e-07 wpdiblcb=-7.846842847e-07 ppdiblcb=1.584128481e-13 drout=1.401076980e+00 ldrout=-1.812387319e-07 wdrout=-1.125811917e-12 pdrout=2.268084520e-19 pscbe1=5.671683714e+09 lpscbe1=-9.852325431e+02 wpscbe1=-4.092825458e+03 ppscbe1=8.262636962e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.181956457e-05 lalpha0=1.046574614e-11 walpha0=4.362788622e-11 palpha0=-8.807641298e-18 alpha1=0.85 beta0=-4.222688583e+01 lbeta0=1.141574186e-05 wbeta0=4.687461261e-05 pbeta0=-9.463093669e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.851246078e-01 lkt1=-1.127225419e-08 wkt1=-9.229597691e-08 pkt1=1.863280410e-14 kt2=-3.744743046e-02 lkt2=1.729815628e-09 wkt2=-4.152799810e-09 pkt2=8.383713756e-16 at=5.963692584e+05 lat=-1.145975016e-01 wat=-4.450171553e-01 pat=8.984050834e-8 ute=-2.073227499e-02 lute=-2.621043079e-07 wute=-9.507226638e-07 pute=1.919328421e-13 ua1=5.505935893e-09 lua1=-1.116358167e-15 wua1=-2.952993833e-15 pua1=5.961533475e-22 ub1=-2.441486443e-18 lub1=6.357716432e-25 wub1=5.395506944e-25 pub1=-1.089250345e-31 uc1=4.003702278e-10 luc1=-5.111303463e-17 wuc1=-3.772222153e-16 puc1=7.615399807e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.79 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.708872316e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.136298490e-09 wvth0=-4.523411464e-08 pvth0=-2.331164699e-14 k1=9.070734929e-01 lk1=-3.812541394e-16 wk1=-2.432173574e-15 pk1=3.207576427e-22 k2=-2.149820887e-01 lk2=2.026419379e-08 wk2=3.810607722e-08 pk2=-1.071865402e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587083017e-01 ldsub=-1.580764761e-11 wdsub=-5.804669759e-11 pdsub=1.171855116e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000029e-03 lcdscd=-4.034331029e-18 wcdscd=-2.446815667e-17 pcdscd=3.394171229e-24 cit=0.0 voff='-1.237493862e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907111e-08 wvoff=9.859357775e-16 pvoff=-1.519409598e-22 nfactor=1.731365944e+01 lnfactor=-2.973153864e-06 wnfactor=-1.122036921e-05 pnfactor=2.265179357e-12 eta0=-9.000623338e-03 leta0=1.957188437e-09 weta0=8.156419615e-09 peta0=-1.646626080e-15 etab=-4.399799988e-02 letab=-1.646163761e-17 wetab=-1.050153298e-16 petab=1.384951875e-23 u0=5.547781049e-02 lu0=-7.217716904e-09 wu0=-1.873112701e-08 pu0=5.343765601e-15 ua=-1.152485641e-09 lua=-4.258349075e-18 wua=-4.156187318e-17 pua=8.390553155e-24 ub=2.691857246e-18 lub=-1.066794211e-25 wub=-4.391850840e-25 pub=8.866312423e-32 uc=-4.041511711e-10 luc=1.002765479e-16 wuc=3.899493811e-16 puc=-7.872337099e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.043255830e+04 lvsat=1.837387422e-02 wvsat=9.230964961e-02 pvsat=-1.268751625e-8 a0=1.500000009e+00 la0=-1.164661256e-15 wa0=-7.429843407e-15 pa0=9.798553080e-22 ags=1.250000002e+00 lags=-2.493649731e-16 wags=-1.590798604e-15 pags=2.097957363e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.275885499e-03 lketa=-1.704357844e-08 wketa=-1.410050188e-07 pketa=2.846623422e-14 dwg=0.0 dwb=0.0 pclm=1.138804918e+00 lpclm=-1.817403256e-07 wpclm=-5.847582668e-07 ppclm=1.180515837e-13 pdiblc1=3.569721485e-01 lpdiblc1=1.993876175e-16 wpdiblc1=1.271972749e-15 ppdiblc1=-1.677491479e-22 pdiblc2=8.406112141e-03 lpdiblc2=-5.346036114e-18 wpdiblc2=-3.410449700e-17 ppdiblc2=4.497735517e-24 pdiblcb=-1.032957699e-01 lpdiblcb=-1.582922682e-17 wpdiblcb=-1.009810013e-16 ppdiblcb=1.331748600e-23 drout=5.033266680e-01 ldrout=-1.056039478e-15 wdrout=-6.736900815e-15 pdrout=8.884692981e-22 pscbe1=7.914198808e+08 lpscbe1=-1.043276787e-07 wpscbe1=-6.655502319e-07 ppscbe1=8.777308464e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.389195394e-07 lalpha0=-2.368458626e-14 walpha0=-9.870350954e-14 palpha0=1.992636348e-20 alpha1=0.85 beta0=1.174327808e+01 lbeta0=5.201911974e-07 wbeta0=2.548267876e-06 pbeta0=-5.144468673e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.104663883e-01 lkt1=-2.634433021e-08 wkt1=-1.097877690e-07 pkt1=2.216406458e-14 kt2=-2.887893895e-02 lkt2=-6.328021440e-18 wkt2=-4.036893042e-17 pkt2=5.323907981e-24 at=-1.293342571e+05 lat=3.190824978e-02 wat=8.225292804e-02 pat=-1.660530336e-8 ute=-1.273184334e+00 lute=-9.258033808e-09 wute=-3.858207308e-08 pute=7.788987519e-15 ua1=-2.384732695e-11 lua1=-1.193990495e-24 wua1=-7.616946105e-24 pua1=1.004530469e-30 ub1=7.077531829e-19 lub1=-1.696121050e-33 wub1=-1.082023958e-32 pub1=1.426983896e-39 uc1=1.471862498e-10 luc1=2.455868219e-26 wuc1=1.566696624e-25 puc1=-2.066173093e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.80 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='1.769632751e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.397673593e-07 wvth0=-9.137795170e-07 pvth0=9.123298922e-14 k1=0.90707349 k2=3.289612822e-03 lk2=-8.521696480e-09 wk2=-1.582013346e-07 pk2=1.517056376e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.584472951e-01 ldsub=1.861415691e-11 wdsub=1.354431545e-10 pdsub=-1.379908403e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999994e-03 lcdscd=6.320942034e-19 wcdscd=5.300850037e-18 pcdscd=-5.317950941e-25 cit=0.0 voff='-2.075299991e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.845946198e-17 wvoff=-7.304885585e-16 pvoff=7.442291228e-23 nfactor=-2.913988266e+01 lnfactor=3.153185722e-06 wnfactor=2.398368113e-05 pnfactor=-2.377566006e-12 eta0=2.567257691e-02 leta0=-2.615547546e-09 weta0=-1.903164350e-08 peta0=1.938962872e-15 etab=-0.043998 u0=-5.173673152e-02 lu0=6.921844110e-09 wu0=7.362145915e-08 pu0=-6.835785814e-15 ua=-7.206724688e-10 lua=-6.120630210e-17 wua=-2.711245794e-16 pua=3.866551242e-23 ub=1.771516367e-18 lub=1.469605428e-26 wub=4.018009124e-25 pub=-2.224694996e-32 uc=1.304381426e-09 luc=-1.250464396e-16 wuc=-9.098818885e-16 puc=9.269967669e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.037410638e+05 lvsat=7.387065213e-03 wvsat=5.892194530e-02 pvsat=-8.284312417e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-4.708175463e-01 lketa=4.521657543e-08 wketa=3.290117110e-07 pketa=-3.352004213e-14 dwg=0.0 dwb=0.0 pclm=-8.890118050e-01 lpclm=8.569017167e-08 wpclm=8.615453093e-07 ppclm=-7.268837818e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.806722828e-07 lalpha0=3.165160284e-14 walpha0=2.303081980e-13 palpha0=-2.346402953e-20 alpha1=0.85 beta0=1.909329699e+01 lbeta0=-4.491366453e-07 wbeta0=-4.132082319e-06 pbeta0=3.665643968e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.365500159e-01 lkt1=1.665990469e-08 wkt1=1.645535608e-07 pkt1=-1.401634433e-14 kt2=-0.028878939 at=3.126140564e+05 lat=-2.637633575e-02 wat=-1.919234987e-01 pat=1.955335797e-8 ute=-2.134844679e+00 lute=1.043785942e-07 wute=5.434938541e-07 pute=-6.897576784e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.81 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.82 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.257996689e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.325072873e-06 wvth0=3.221288904e-08 pvth0=-6.427077288e-13 k1=7.639711556e-01 lk1=-3.909839147e-06 wk1=-9.885369208e-08 pk1=1.972317101e-12 k2=-1.383209333e-01 lk2=1.967761991e-06 wk2=5.361042226e-08 pk2=-1.069628765e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.386994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.069675642e-07 wvoff=2.409444893e-08 pvoff=-4.807295779e-13 nfactor=2.191954229e+00 lnfactor=1.377968224e-05 wnfactor=6.077045009e-07 pnfactor=-1.212484788e-11 eta0=0.08 etab=-0.07 u0=2.273004585e-02 lu0=7.823639617e-08 wu0=1.444533578e-09 pu0=-2.882116205e-14 ua=-1.850827749e-09 lua=1.583145143e-14 wua=3.944440551e-16 pua=-7.869900849e-21 ub=2.674812262e-18 lub=-1.739525219e-23 wub=-4.923778716e-25 pub=9.823864701e-30 uc=6.609339935e-11 luc=-3.502831907e-16 wuc=-1.845083865e-18 puc=3.681289372e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.202541567e+00 la0=3.193466813e-06 wa0=1.226358632e-07 pa0=-2.446816150e-12 ags=5.084562099e-01 lags=-3.263653074e-06 wags=-1.221345977e-07 pags=2.436814959e-12 a1=0.0 a2=0.42385546 b0=3.944133822e-07 lb0=-6.602962931e-12 wb0=-2.141577111e-13 pb0=4.272849167e-18 b1=1.182299395e-08 lb1=-1.856241993e-13 wb1=-5.659323710e-15 pb1=1.129141532e-19 keta=-3.460253357e-02 lketa=5.996724100e-07 wketa=2.080089353e-08 pketa=-4.150169524e-13 dwg=0.0 dwb=0.0 pclm=-1.551262420e-01 lpclm=3.431748312e-06 wpclm=9.476407614e-08 ppclm=-1.890721570e-12 pdiblc1=0.39 pdiblc2=-8.044955951e-03 lpdiblc2=1.796723430e-07 wpdiblc2=5.599972445e-09 ppdiblc2=-1.117299838e-13 pdiblcb=1.194793931e+01 lpdiblcb=-2.388826604e-04 wpdiblcb=-7.798238780e-06 ppdiblcb=1.555895322e-10 drout=0.56 pscbe1=-5.454128204e+08 lpscbe1=1.537118491e+04 wpscbe1=3.075658461e+02 ppscbe1=-6.136517161e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.759117059e-01 lkt1=-2.088621580e-07 wkt1=-4.763800346e-09 pkt1=9.504677761e-14 kt2=-3.508984941e-02 lkt2=1.111702531e-07 wkt2=-2.322708176e-10 pkt2=4.634239713e-15 at=1.981929863e+05 lat=-4.627437017e-1 ute=-8.928439532e-01 lute=-4.440411761e-06 wute=-8.034469240e-08 pute=1.603027742e-12 ua1=5.088873862e-10 lua1=1.221279803e-14 wua1=3.395096515e-16 pua1=-6.773856166e-21 ub1=1.164653596e-19 lub1=-1.368570067e-23 wub1=-3.254671057e-25 pub1=6.493680963e-30 uc1=9.556390960e-11 luc1=-1.231939818e-15 wuc1=-1.716993806e-17 puc1=3.425725610e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.83 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.902240806e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.758951840e-08 wvth0=-4.784370729e-08 pvth0=-6.107201538e-15 k1=5.991074590e-01 lk1=-2.598862650e-06 wk1=-1.053621493e-07 pk1=2.024071578e-12 k2=-9.734850519e-03 lk2=9.452607626e-07 wk2=1.315076145e-08 pk2=-7.478983572e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077859692e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.611475537e-07 wvoff=-6.652270698e-09 pvoff=-2.362353222e-13 nfactor=6.691706598e+00 lnfactor=-2.200181313e-05 wnfactor=-3.086819217e-06 pnfactor=1.725356507e-11 eta0=0.08 etab=-0.07 u0=5.016141404e-02 lu0=-1.398945793e-07 wu0=-1.457667305e-08 pu0=9.857756652e-14 ua=1.921968839e-09 lua=-1.416937807e-14 wua=-1.889104298e-15 pua=1.028860392e-20 ub=-7.838765265e-19 lub=1.010782947e-23 wub=1.682484813e-24 pub=-7.470384556e-30 uc=1.457305801e-10 luc=-9.835485750e-16 wuc=-8.859884428e-17 puc=7.266684729e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.030118304e+00 la0=-3.387324923e-06 wa0=-4.046018659e-07 pa0=1.745715531e-12 ags=2.965423767e-01 lags=-1.578539491e-06 wags=4.204292826e-08 pags=1.131294810e-12 a1=0.0 a2=0.42385546 b0=-1.899679869e-07 lb0=-1.956031826e-12 wb0=1.408274480e-13 pb0=1.450049425e-18 b1=5.717141510e-09 lb1=-1.370711873e-13 wb1=-4.238242778e-15 pb1=1.016138867e-19 keta=2.140568848e-02 lketa=1.543016932e-07 wketa=-2.527657375e-08 pketa=-4.861441587e-14 dwg=0.0 dwb=0.0 pclm=2.022332362e+00 lpclm=-1.388314339e-05 wpclm=-1.766586218e-06 ppclm=1.291051447e-11 pdiblc1=0.39 pdiblc2=3.611915776e-02 lpdiblc2=-1.715154337e-07 wpdiblc2=-2.458276908e-08 ppdiblc2=1.282795851e-13 pdiblcb=-3.594381794e+01 lpdiblcb=1.419468942e-04 wpdiblcb=2.339471634e-05 ppdiblcb=-9.245313501e-11 drout=0.56 pscbe1=1.778990503e+09 lpscbe1=-3.112193713e+03 wpscbe1=-7.423504445e+02 ppscbe1=2.212292242e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.272022175e-01 lkt1=1.989938870e-07 wkt1=2.664120078e-08 pkt1=-1.546820541e-13 kt2=-9.811760398e-02 lkt2=6.123594571e-07 wkt2=5.748353971e-08 pkt2=-4.543150175e-13 at=140000.0 ute=-3.341961982e+00 lute=1.503468336e-05 wute=1.374777495e-06 pute=-9.967930737e-12 ua1=-6.388335101e-10 lua1=2.133933802e-14 wua1=1.402402819e-15 pua1=-1.522585615e-20 ub1=-2.813180195e-19 lub1=-1.052257457e-23 wub1=-4.852743371e-25 pub1=7.764449050e-30 uc1=2.621286344e-10 luc1=-2.556442688e-15 wuc1=-2.169010355e-16 puc1=1.930810480e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.84 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='3.582951813e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.341449290e-07 wvth0=1.116558878e-07 pvth0=-6.364306210e-13 k1=-4.042235728e-01 lk1=1.366182191e-06 wk1=6.275222338e-07 pk1=-8.722002908e-13 k2=3.812518825e-01 lk2=-5.998722788e-07 wk2=-2.715107787e-07 pk2=3.770501747e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.558838394e+00 ldsub=8.373397193e-06 wdsub=1.570741516e-06 pdsub=-6.207383554e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.777900094e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.162602830e-06 wvoff=-2.701670131e-07 pvoff=8.051435816e-13 nfactor=5.659190481e+00 lnfactor=-1.792143230e-05 wnfactor=-1.773617076e-06 pnfactor=1.206394648e-11 eta0=-4.814921745e-01 leta0=2.218950256e-06 weta0=4.162465018e-07 peta0=-1.644956642e-12 etab=4.208642281e-01 letab=-1.939837016e-06 wetab=-3.638884513e-07 petab=1.438043857e-12 u0=2.034160379e-02 lu0=-2.205023777e-08 wu0=6.919807228e-09 pu0=1.362603455e-14 ua=3.029379355e-09 lua=-1.854573265e-14 wua=-2.432595795e-15 pua=1.243641763e-20 ub=-5.138495807e-18 lub=2.731676667e-23 wub=4.498493139e-24 pub=-1.859891436e-29 uc=-2.799473311e-10 luc=6.986798745e-16 wuc=2.055672917e-16 puc=-4.358410906e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=-3.638847673e-01 la0=6.073490330e-06 wa0=1.282985179e-06 pa0=-4.923427648e-12 ags=-6.469315077e-01 lags=2.149957027e-06 wags=6.347997239e-07 pags=-1.211209509e-12 a1=0.0 a2=0.42385546 b0=-3.646607291e-07 lb0=-1.265666897e-12 wb0=2.703310210e-13 pb0=9.382667155e-19 b1=3.314007703e-09 lb1=-1.275742885e-13 wb1=-2.456746818e-15 pb1=9.457362670e-20 keta=2.259918777e-01 lketa=-6.541985807e-07 wketa=-1.468382588e-07 pketa=4.317828977e-13 dwg=0.0 dwb=0.0 pclm=-3.852630753e+00 lpclm=9.334011723e-06 wpclm=3.233970149e-06 ppclm=-6.851089229e-12 pdiblc1=0.39 pdiblc2=-6.257524983e-03 lpdiblc2=-4.047826320e-09 wpdiblc2=5.705853750e-09 ppdiblc2=8.582551968e-15 pdiblcb=6.328493310e-02 lpdiblcb=-3.488915497e-07 wpdiblcb=-6.544756318e-08 ppdiblcb=2.586409814e-13 drout=0.56 pscbe1=1.178330128e+09 lpscbe1=-7.384553890e+02 wpscbe1=-3.606941876e+02 ppscbe1=7.040321316e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-5.599990113e-01 lkt1=1.118979113e-06 wkt1=1.959372255e-07 pkt1=-8.237197976e-13 kt2=-8.630210486e-02 lkt2=5.656660106e-07 wkt2=4.646331980e-08 pkt2=-4.107644198e-13 at=1.551821722e+05 lat=-5.999813783e-02 wat=9.581523249e-03 pat=-3.786503968e-8 ute=-7.911511772e+00 lute=3.309300035e-05 wute=4.580579668e-06 pute=-2.263687943e-11 ua1=-2.072426389e-08 lua1=1.007145687e-13 wua1=1.488308955e-14 pua1=-6.849992591e-20 ub1=1.724441975e-17 lub1=-7.978220469e-23 wub1=-1.219309854e-23 pub1=5.403237706e-29 uc1=-1.177121865e-10 luc1=-1.055356965e-15 wuc1=8.234223907e-17 puc1=7.482366687e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.85 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='8.144787272e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.372893329e-08 wvth0=-2.167794065e-07 pvth0=4.635989689e-15 k1=6.370895852e-01 lk1=-6.663371774e-07 wk1=-2.995472631e-08 pk1=4.111164956e-13 k2=-8.267798593e-03 lk2=1.604237858e-07 wk2=-3.089019493e-08 pk2=-9.261257094e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.083241089e+00 ldsub=-4.591151551e-06 wdsub=-3.141483033e-06 pdsub=2.990318010e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.614723649e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.516125218e-08 wvoff=1.926616597e-07 pvoff=-9.824291114e-14 nfactor=-3.850612951e-01 lnfactor=-6.123772104e-06 wnfactor=2.391445590e-06 pnfactor=3.934239800e-12 eta0=1.276724988e+00 leta0=-1.212880418e-06 weta0=-8.324927483e-07 peta0=7.924337744e-13 etab=-1.038045167e+00 letab=9.077805120e-07 wetab=7.277769025e-07 petab=-6.927570058e-13 u0=7.455837770e-03 lu0=3.101244091e-09 wu0=1.635482177e-08 pu0=-4.789991066e-15 ua=-9.544789026e-09 lua=5.997547707e-15 wua=6.383127579e-15 pua=-4.770825321e-21 ub=1.384985332e-17 lub=-9.746231213e-24 wub=-8.817880785e-24 pub=7.393062895e-30 uc=-1.252442974e-10 luc=3.967179623e-16 wuc=1.216217375e-16 puc=-2.719893585e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.512613283e+04 lvsat=1.071072587e-01 wvsat=3.362270169e-02 pvsat=-6.562751260e-8 a0=7.974719482e+00 la0=-1.020247287e-05 wa0=-4.864090681e-06 pa0=7.074932929e-12 ags=4.395513928e+00 lags=-7.692296413e-06 wags=-3.032158887e-06 pags=5.946257332e-12 a1=0.0 a2=0.42385546 b0=-6.430353943e-07 lb0=-7.223126771e-13 wb0=4.766962846e-13 pb0=5.354662784e-19 b1=-7.787721762e-08 lb1=3.090132157e-14 wb1=5.773209472e-14 pb1=-2.290782951e-20 keta=-7.196537533e-01 lketa=1.191589159e-06 wketa=5.139678209e-07 pketa=-8.580319340e-13 dwg=0.0 dwb=0.0 pclm=2.412891835e+00 lpclm=-2.895542771e-06 wpclm=-1.468342163e-06 ppclm=2.327264830e-12 pdiblc1=5.467295616e-01 lpdiblc1=-3.059174535e-07 wpdiblc1=-7.999047045e-08 ppdiblc1=1.561318794e-13 pdiblc2=-2.944953112e-02 lpdiblc2=4.122020981e-08 wpdiblc2=2.539859168e-08 ppdiblc2=-2.985532904e-14 pdiblcb=1.604222365e-01 lpdiblcb=-5.384920065e-07 wpdiblcb=-1.202590924e-07 ppdiblcb=3.656265638e-13 drout=4.313542261e+00 ldrout=-7.326467821e-06 wdrout=-2.667774013e-06 pdrout=5.207177409e-12 pscbe1=3.446387392e+08 lpscbe1=8.888109931e+02 wpscbe1=3.375693206e+02 ppscbe1=-6.588951430e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.785825191e-05 lalpha0=-7.383624616e-11 walpha0=-2.804206858e-11 palpha0=5.473478086e-17 alpha1=2.049605555e+00 lalpha1=-2.341487291e-06 walpha1=-7.813294895e-07 palpha1=1.525062185e-12 beta0=3.868679618e+01 lbeta0=-4.845895175e-05 wbeta0=-1.840465020e-05 pbeta0=3.592368703e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=1.461049701e-01 lkt1=-2.592518322e-07 wkt1=-3.492656170e-07 pkt1=2.404512719e-13 kt2=4.943918352e-01 lkt2=-5.677794577e-07 wkt2=-3.665497230e-07 pkt2=3.953878913e-13 at=2.683129784e+03 lat=2.376618456e-01 wat=9.842944184e-02 pat=-2.112856039e-7 ute=1.845552780e+01 lute=-1.837232321e-05 wute=-1.355411642e-05 pute=1.275988930e-11 ua1=5.931986210e-08 lua1=-5.552203995e-14 wua1=-3.962998783e-14 pua1=3.790311408e-20 ub1=-4.472169872e-17 lub1=4.116828460e-23 wub1=2.973571533e-23 pub1=-2.780767808e-29 uc1=-1.144071374e-09 luc1=9.479740314e-16 wuc1=7.916638482e-16 puc1=-6.362747030e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.86 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='1.150217030e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.758539786e-07 wvth0=-4.034244171e-07 pvth0=1.822998290e-13 k1=-5.490799469e-01 lk1=4.627550630e-07 wk1=7.652063214e-07 pk1=-3.457821977e-13 k2=3.166869134e-01 lk2=-1.488944304e-07 wk2=-2.440327212e-07 pk2=1.102737501e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790972e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.880217007e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.104330605e-07 wvoff=1.702961243e-07 pvoff=-7.695358295e-14 nfactor=-1.563230129e+01 lnfactor=8.389785953e-06 wnfactor=1.242122284e-05 pnfactor=-5.612914598e-12 eta0=-4.380236984e-01 leta0=4.193562769e-07 weta0=-5.106728688e-13 peta0=2.307633667e-19 etab=-1.600650675e-01 letab=7.204793715e-8 u0=-2.204651287e-03 lu0=1.229688008e-08 wu0=2.155570607e-08 pu0=-9.740614014e-15 ua=-4.867405384e-09 lua=1.545235089e-15 wua=2.610305085e-15 pua=-1.179547272e-21 ub=4.976298969e-18 lub=-1.299663426e-24 wub=-2.001020570e-24 pub=9.042231761e-31 uc=5.075196463e-10 luc=-2.055980132e-16 wuc=-3.124398747e-16 puc=1.411856430e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.263343699e+05 lvsat=1.076906086e-02 wvsat=-6.724540339e-02 pvsat=3.038692013e-8 a0=-6.474326697e+00 la0=3.551299655e-06 wa0=4.889794855e-06 pa0=-2.209605389e-12 ags=-7.157793252e+00 lags=3.305077179e-06 wags=6.120005796e-06 pags=-2.765514339e-12 a1=0.0 a2=0.42385546 b0=-2.668811703e-06 lb0=1.205985301e-12 wb0=1.978448829e-12 pb0=-8.940234353e-19 b1=-8.645704443e-08 lb1=3.906829570e-14 wb1=6.409250909e-14 pb1=-2.896218710e-20 keta=1.019557592e+00 lketa=-4.639330751e-07 wketa=-7.375914614e-07 pketa=3.333035671e-13 dwg=0.0 dwb=0.0 pclm=-1.605842467e+00 lpclm=9.298140543e-07 wpclm=1.859155647e-06 ppclm=-8.401171128e-13 pdiblc1=3.991551774e-01 lpdiblc1=-1.654442010e-07 wpdiblc1=1.599809409e-07 ppdiblc1=-7.229234755e-14 pdiblc2=2.633355276e-02 lpdiblc2=-1.187864786e-08 wpdiblc2=-1.135778438e-08 ppdiblc2=5.132366963e-15 pdiblcb=-6.860776615e-01 lpdiblcb=2.672751629e-07 wpdiblcb=5.023084374e-07 ppdiblcb=-2.269836390e-13 drout=-7.344739711e+00 ldrout=3.770829280e-06 wdrout=5.335548027e-06 pdrout=-2.411032778e-12 pscbe1=2.038836018e+09 lpscbe1=-7.238632065e+02 wpscbe1=-6.751386411e+02 ppscbe1=3.050823243e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-7.912406276e-05 lalpha0=3.751699650e-11 walpha0=5.608413716e-11 palpha0=-2.534335598e-17 alpha1=-1.549211111e+00 lalpha1=1.084157916e-06 walpha1=1.562658979e-06 palpha1=-7.061359021e-13 beta0=-3.955143475e+01 lbeta0=2.601453375e-05 wbeta0=3.680930040e-05 pbeta0=-1.663342347e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=1.174945592e-02 lkt1=-1.313613710e-07 wkt1=-1.840160659e-07 pkt1=8.315336386e-14 kt2=-1.611696512e-01 lkt2=5.623706546e-08 wkt2=9.295234878e-08 pkt2=-4.200340032e-14 at=4.708019125e+05 lat=-2.079315295e-01 wat=-2.351849767e-01 pat=1.062756224e-7 ute=-4.255336348e-01 lute=-3.997995752e-07 wute=-2.840331857e-07 pute=1.283492000e-13 ua1=1.135188042e-09 lua1=-1.371542308e-16 wua1=3.601632756e-16 pua1=-1.627509412e-22 ub1=-2.231833164e-18 lub1=7.229888876e-25 wub1=9.943687287e-25 pub1=-4.493363355e-31 uc1=-2.872795245e-10 luc1=1.324101492e-16 wuc1=2.345901449e-16 puc1=-1.060068293e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.87 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.883840693e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.197233829e-8 k1=1.260614571e-01 lk1=1.576714902e-7 k2=8.571419420e-02 lk2=-4.452224711e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458427e-8 nfactor=3.214803974e+00 lnfactor=-1.268628226e-7 eta0=8.851262253e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 wetab=9.540979118e-24 petab=1.301042607e-30 u0=2.084392174e-02 lu0=1.881667846e-9 ua=-1.669318486e-09 lua=1.000803833e-16 ub=2.049104468e-18 lub=2.308015275e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.493390954e+05 lvsat=3.736624816e-4 a0=1.291411731e+00 la0=4.211000822e-8 ags=-7.269793732e-01 lags=3.991145728e-07 pags=5.551115123e-29 a1=0.0 a2=0.42385546 b0=-1.068120851e-16 lb0=2.156333055e-23 b1=2.864312598e-18 lb1=-5.782502915e-25 keta=5.428652146e-02 lketa=-2.774541862e-08 wketa=2.775557562e-23 pketa=8.673617380e-30 dwg=0.0 dwb=0.0 pclm=6.240064173e-01 lpclm=-7.781228934e-8 pdiblc1=-2.285578198e-01 lpdiblc1=1.182073759e-07 wpdiblc1=5.551115123e-23 ppdiblc1=2.775557562e-29 pdiblc2=-6.704200072e-03 lpdiblc2=3.050484931e-09 wpdiblc2=-2.222614454e-24 ppdiblc2=1.599198204e-30 pdiblcb=-8.758737421e-02 lpdiblcb=-3.171226653e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016608e+08 lpscbe1=1.293488348e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901082e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-9 at=-3.932844299e+03 lat=6.592087176e-03 pat=3.637978807e-24 ute=-1.303201518e+00 lute=-3.198134688e-9 ua1=1.522520005e-09 lua1=-3.121821852e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 pub1=1.925929944e-46 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=3.877409121e-32 puc1=-1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.88 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142908321e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442070405e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220557072e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571054398e-16 ags=1.250000000e+00 lags=3.363842538e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689626299e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211488351e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135236432e-18 drout=5.033266589e-01 ldrout=1.424533824e-16 pscbe1=7.914198799e+08 lpscbe1=1.407337189e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.536088503e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610623275e-25 ub1=7.077531683e-19 lub1=2.287970107e-34 uc1=1.471862500e-10 luc1=-3.312806654e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.89 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-5.295351531e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.239560175e-07 wvth0=7.906442316e-07 pvth0=-1.042709519e-13 k1=0.90707349 k2=-3.448034743e-01 lk2=2.970539255e-08 wk2=9.984772892e-08 pk2=-1.316801834e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999998e-03 lcdscd=2.454347489e-19 wcdscd=1.858915799e-18 pcdscd=-2.451563258e-25 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193267707e-17 nfactor=6.176567708e+00 lnfactor=-4.448895625e-07 wnfactor=-2.197180485e-06 pnfactor=2.897663596e-13 eta0=8.801660331e-10 leta0=-8.964943129e-17 weta0=4.866420979e-19 peta0=-6.417884652e-26 etab=-0.043998 u0=1.790423397e-01 lu0=-1.963736632e-08 wu0=-9.746014345e-08 pu0=1.285314118e-14 ua=-5.898554346e-10 lua=-7.453406508e-17 wua=-3.681021249e-16 pua=4.854567633e-23 ub=3.153859100e-18 lub=-1.261382387e-25 wub=-6.229601672e-25 pub=8.215660981e-32 uc=7.700399988e-11 luc=1.171427334e-26 wuc=-1.275926095e-28 puc=1.685380498e-35 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.818455598e+05 lvsat=-3.606287063e-03 wvsat=1.021364113e-03 pvsat=-1.346985206e-10 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000006e-02 lketa=6.295533539e-18 wketa=7.294165272e-20 pketa=-9.603429163e-27 dwg=0.0 dwb=0.0 pclm=9.515324736e-01 lpclm=-1.018263203e-07 wpclm=-5.028906565e-07 ppclm=6.632172266e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.406312920e-24 walpha0=-1.457955460e-25 palpha0=1.921705999e-32 alpha1=0.85 beta0=1.103149680e+01 lbeta0=3.734391265e-07 wbeta0=1.844307516e-06 pbeta0=-2.432291195e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-9.125600823e-02 lkt1=-1.851100502e-08 wkt1=-9.142048357e-08 pkt1=1.205662479e-14 kt2=-0.028878939 at=5.372048693e+04 lat=6.909715012e-12 wat=-3.096647561e-14 pat=4.103640094e-21 ute=-2.023669003e+00 lute=9.335978203e-08 wute=4.610768797e-07 pute=-6.080727997e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.90 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.91 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-08 wu0=-2.220446049e-22 ua=-1.245222449e-09 lua=3.748486558e-15 ub=1.918845364e-18 lub=-2.312290614e-24 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-07 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+03 ppscbe1=-1.525878906e-17 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.92 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-07 pk2=-8.881784197e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917323e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 keta=-1.740241834e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 wpclm=-8.881784197e-22 ppclm=1.065814104e-26 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-08 ppdiblc2=-1.110223025e-28 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.93 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872697e-01 leta0=-3.066156572e-7 etab=-1.378278647e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-06 wa0=-1.421085472e-20 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312433e-10 lb1=1.762827905e-14 keta=5.453875497e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-1 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 ub1=-1.476118686e-18 lub1=3.175805416e-24 pub1=1.232595164e-44 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.94 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-09 peta0=6.938893904e-30 etab=7.933901887e-02 letab=-1.558362640e-07 wetab=-1.387778781e-22 petab=2.151057110e-28 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775476e-01 lags=1.437223750e-6 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 keta=6.946103312e-02 lketa=-1.257806426e-07 wketa=1.665334537e-22 pketa=1.665334537e-28 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=2.117582368e-27 palpha0=-4.658681210e-33 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-6 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=1.654361225e-30 pua1=-4.963083675e-36 ub1=9.327016030e-19 lub1=-1.525925138e-24 wub1=-3.081487911e-39 pub1=3.081487911e-45 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.95 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.308238316e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.038039511e-9 k1=6.257710814e-01 lk1=-6.813779454e-8 k2=-5.798601513e-02 lk2=2.041314719e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790972e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594373e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716768537e-9 nfactor=3.438485258e+00 lnfactor=-2.279401452e-7 eta0=-4.380244825e-01 leta0=4.193566312e-07 peta0=-1.360023205e-27 etab=-1.600650675e-01 letab=7.204793715e-8 u0=3.089066266e-02 lu0=-2.658263485e-9 ua=-8.597024590e-10 lua=-2.657697166e-16 ub=1.904054258e-18 lub=8.862558670e-26 uc=2.781855420e-11 luc=1.116979601e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.308988651e+04 lvsat=5.742328124e-2 a0=1.033165535e+00 la0=1.588065578e-7 ags=2.238489687e+00 lags=-9.409245514e-7 a1=0.0 a2=0.42385546 b0=3.687777371e-07 lb0=-1.666436526e-13 b1=1.194667768e-08 lb1=-5.398476655e-15 keta=-1.128952678e-01 lketa=4.780085550e-8 dwg=0.0 dwb=0.0 pclm=1.248591510e+00 lpclm=-3.600504257e-7 pdiblc1=6.447801384e-01 lpdiblc1=-2.764374541e-7 pdiblc2=8.895504641e-03 lpdiblc2=-3.998725234e-9 pdiblcb=8.513601992e-02 lpdiblcb=-8.122164671e-08 wpdiblcb=-1.196959198e-22 ppdiblcb=8.326672685e-29 drout=8.471347030e-01 ldrout=6.907687805e-8 pscbe1=1.002269402e+09 lpscbe1=-2.554584477e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094440e-06 lalpha0=-1.393643679e-12 alpha1=0.85 beta0=1.696331585e+01 lbeta0=4.765917258e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775674e-01 lkt1=-3.692777228e-9 kt2=-1.845629469e-02 lkt2=-8.252388786e-9 at=1.097132702e+05 lat=-4.476243271e-2 ute=-8.616208324e-01 lute=-2.027400563e-7 ua1=1.688160728e-09 lua1=-3.870320810e-16 wua1=1.323488980e-29 ub1=-7.051401785e-19 lub1=3.310533463e-26 uc1=7.289584949e-11 luc1=-3.034625898e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.96 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.883840693e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.197233829e-8 k1=1.260614571e-01 lk1=1.576714902e-7 k2=8.571419420e-02 lk2=-4.452224711e-08 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458427e-8 nfactor=3.214803974e+00 lnfactor=-1.268628226e-07 wnfactor=-2.842170943e-20 eta0=8.851262253e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 wetab=-1.387778781e-23 petab=5.204170428e-29 u0=2.084392174e-02 lu0=1.881667846e-9 ua=-1.669318486e-09 lua=1.000803833e-16 ub=2.049104468e-18 lub=2.308015275e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.493390954e+05 lvsat=3.736624816e-4 a0=1.291411731e+00 la0=4.211000822e-8 ags=-7.269793732e-01 lags=3.991145728e-07 pags=1.332267630e-27 a1=0.0 a2=0.42385546 b0=-1.068120851e-16 lb0=2.156333055e-23 b1=2.864312598e-18 lb1=-5.782502915e-25 keta=5.428652146e-02 lketa=-2.774541862e-08 wketa=-1.110223025e-22 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=6.240064173e-01 lpclm=-7.781228934e-8 pdiblc1=-2.285578198e-01 lpdiblc1=1.182073759e-07 wpdiblc1=-4.440892099e-22 ppdiblc1=1.110223025e-28 pdiblc2=-6.704200072e-03 lpdiblc2=3.050484931e-09 wpdiblc2=-1.517883041e-23 ppdiblc2=1.626303259e-30 pdiblcb=-8.758737421e-02 lpdiblcb=-3.171226653e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016608e+08 lpscbe1=1.293488348e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901082e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-9 at=-3.932844299e+03 lat=6.592087176e-3 ute=-1.303201518e+00 lute=-3.198134688e-9 ua1=1.522520005e-09 lua1=-3.121821852e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 pub1=1.540743956e-45 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=-2.067951531e-31 puc1=3.877409121e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.97 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.143263593e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442105100e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220446049e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571081043e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689581891e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211453656e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135180921e-18 drout=5.033266589e-01 ldrout=1.424531604e-16 pscbe1=7.914198799e+08 lpscbe1=1.407241821e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.535394613e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610624050e-25 ub1=7.077531683e-19 lub1=2.287973959e-34 uc1=1.471862500e-10 luc1=-3.312444763e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.98 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='9.297747778e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.172075883e-06 wvth0=-5.610081341e-06 pvth0=7.398631374e-13 k1=0.90707349 k2=5.762027147e-01 lk2=-9.175782466e-08 wk2=-5.000238641e-07 pk2=6.594364722e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000021e-03 lcdscd=-2.688169132e-18 wcdscd=-1.262934202e-17 pcdscd=1.665570459e-24 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193356525e-17 nfactor=6.176568640e+00 lnfactor=-4.448896854e-07 wnfactor=-2.197181092e-06 pnfactor=2.897664396e-13 eta0=8.801661157e-10 leta0=-8.964943057e-17 weta0=4.866456862e-19 peta0=-6.417931974e-26 etab=-0.043998 u0=-8.366923922e-01 lu0=1.143187459e-07 wu0=5.641102336e-07 pu0=-7.439542171e-14 ua=-5.898507852e-10 lua=-7.453467825e-17 wua=-3.681051531e-16 pua=4.854607570e-23 ub=3.153933276e-18 lub=-1.261480212e-25 wub=-6.230084797e-25 pub=8.216298132e-32 uc=7.700399988e-11 luc=1.191553672e-26 wuc=8.652309207e-28 puc=-1.141509245e-34 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-8.301504799e+05 lvsat=1.298567626e-01 wvsat=6.601566487e-01 pvsat=-8.706211898e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000006e-02 lketa=6.180167489e-18 wketa=-4.964917366e-19 pketa=6.550315845e-26 dwg=0.0 dwb=0.0 pclm=9.515324590e-01 lpclm=-1.018263184e-07 wpclm=-5.028906469e-07 ppclm=6.632172140e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.175575852e-24 walpha0=9.927226142e-25 palpha0=-1.309724695e-31 alpha1=0.85 beta0=1.100264470e+01 lbeta0=3.772441712e-07 wbeta0=1.863099528e-06 pbeta0=-2.457074288e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-8.859297576e-02 lkt1=-1.886220840e-08 wkt1=-9.315497521e-08 pkt1=1.228537129e-14 kt2=-0.028878939 at=5.372048693e+04 lat=6.959075108e-12 wat=2.123415470e-13 pat=-2.805609256e-20 ute=-2.030882020e+00 lute=9.431104186e-08 wute=4.657748760e-07 pute=-6.142685643e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.99 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.100 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-8 ua=-1.245222449e-09 lua=3.748486558e-15 ub=1.918845364e-18 lub=-2.312290614e-24 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-7 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+03 ppscbe1=7.629394531e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.101 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-07 pk2=2.220446049e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917323e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 pb1=2.646977960e-35 keta=-1.740241833e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 wpclm=6.661338148e-22 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 wuc1=1.033975766e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.102 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872697e-01 leta0=-3.066156572e-7 etab=-1.378278648e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-6 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312434e-10 lb1=1.762827905e-14 keta=5.453875497e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-1 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 ub1=-1.476118686e-18 lub1=3.175805416e-24 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.103 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-09 weta0=1.734723476e-24 peta0=1.734723476e-30 etab=7.933901887e-02 letab=-1.558362640e-07 wetab=-6.418476861e-23 petab=5.204170428e-30 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 pua=1.654361225e-36 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775476e-01 lags=1.437223750e-06 pags=1.776356839e-27 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 keta=6.946103312e-02 lketa=-1.257806426e-07 wketa=-2.775557562e-23 pketa=-1.110223025e-28 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=5.505714157e-27 palpha0=-1.694065895e-33 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-6 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=8.271806126e-31 pua1=-1.654361225e-36 ub1=9.327016030e-19 lub1=-1.525925138e-24 wub1=-7.703719778e-40 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.104 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.308238316e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.038039511e-9 k1=6.257710814e-01 lk1=-6.813779454e-08 wk1=-1.776356839e-21 k2=-5.798601513e-02 lk2=2.041314719e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790972e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594373e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716768537e-9 nfactor=3.438485258e+00 lnfactor=-2.279401452e-7 eta0=-4.380244825e-01 leta0=4.193566312e-07 weta0=4.163336342e-23 peta0=3.851086117e-28 etab=-1.600650675e-01 letab=7.204793715e-8 u0=3.089066266e-02 lu0=-2.658263485e-9 ua=-8.597024590e-10 lua=-2.657697166e-16 ub=1.904054258e-18 lub=8.862558670e-26 uc=2.781855420e-11 luc=1.116979601e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.308988651e+04 lvsat=5.742328124e-2 a0=1.033165535e+00 la0=1.588065578e-7 ags=2.238489687e+00 lags=-9.409245514e-7 a1=0.0 a2=0.42385546 b0=3.687777371e-07 lb0=-1.666436526e-13 b1=1.194667768e-08 lb1=-5.398476655e-15 keta=-1.128952678e-01 lketa=4.780085550e-08 pketa=1.110223025e-28 dwg=0.0 dwb=0.0 pclm=1.248591510e+00 lpclm=-3.600504257e-7 pdiblc1=6.447801384e-01 lpdiblc1=-2.764374541e-07 wpdiblc1=1.776356839e-21 pdiblc2=8.895504641e-03 lpdiblc2=-3.998725234e-9 pdiblcb=8.513601992e-02 lpdiblcb=-8.122164671e-08 wpdiblcb=-3.122502257e-23 ppdiblcb=-8.283304598e-29 drout=8.471347030e-01 ldrout=6.907687805e-8 pscbe1=1.002269402e+09 lpscbe1=-2.554584477e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094440e-06 lalpha0=-1.393643679e-12 alpha1=0.85 beta0=1.696331585e+01 lbeta0=4.765917258e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775674e-01 lkt1=-3.692777228e-9 kt2=-1.845629469e-02 lkt2=-8.252388786e-9 at=1.097132702e+05 lat=-4.476243271e-2 ute=-8.616208324e-01 lute=-2.027400563e-7 ua1=1.688160728e-09 lua1=-3.870320810e-16 ub1=-7.051401785e-19 lub1=3.310533463e-26 uc1=7.289584949e-11 luc1=-3.034625898e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.105 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.883840693e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.197233829e-8 k1=1.260614571e-01 lk1=1.576714902e-7 k2=8.571419420e-02 lk2=-4.452224711e-08 wk2=5.551115123e-23 pk2=-4.163336342e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-09 pcdscd=3.469446952e-30 cit=0.0 voff='-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458427e-8 nfactor=3.214803974e+00 lnfactor=-1.268628226e-7 eta0=8.851262253e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 wetab=2.602085214e-23 petab=-1.301042607e-29 u0=2.084392174e-02 lu0=1.881667846e-9 ua=-1.669318486e-09 lua=1.000803833e-16 ub=2.049104468e-18 lub=2.308015275e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.493390954e+05 lvsat=3.736624816e-4 a0=1.291411731e+00 la0=4.211000822e-8 ags=-7.269793732e-01 lags=3.991145728e-07 wags=4.440892099e-22 pags=-1.110223025e-28 a1=0.0 a2=0.42385546 b0=-1.068120851e-16 lb0=2.156333055e-23 b1=2.864312598e-18 lb1=-5.782502915e-25 keta=5.428652146e-02 lketa=-2.774541862e-08 wketa=-2.775557562e-23 pketa=-2.081668171e-29 dwg=0.0 dwb=0.0 pclm=6.240064173e-01 lpclm=-7.781228934e-8 pdiblc1=-2.285578198e-01 lpdiblc1=1.182073759e-07 wpdiblc1=1.110223025e-22 ppdiblc1=8.326672685e-29 pdiblc2=-6.704200072e-03 lpdiblc2=3.050484931e-09 wpdiblc2=-5.204170428e-24 ppdiblc2=1.490777987e-30 pdiblcb=-8.758737421e-02 lpdiblcb=-3.171226653e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016608e+08 lpscbe1=1.293488348e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901082e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-06 wbeta0=5.684341886e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-9 at=-3.932844299e+03 lat=6.592087176e-3 ute=-1.303201518e+00 lute=-3.198134688e-9 ua1=1.522520005e-09 lua1=-3.121821852e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=5.169878828e-32 puc1=-3.231174268e-39 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.106 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142819504e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442070405e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220557072e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571063279e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-08 pketa=-5.551115123e-29 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689626299e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211453656e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135402966e-18 drout=5.033266589e-01 ldrout=1.424531604e-16 pscbe1=7.914198799e+08 lpscbe1=1.407337189e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.535949725e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610623533e-25 ub1=7.077531683e-19 lub1=2.287973959e-34 uc1=1.471862500e-10 luc1=-3.312858353e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.107 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-2.939912633e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.418390099e-07 wvth0=2.238199509e-06 pvth0=-2.951759894e-13 k1=0.90707349 k2=-5.071645056e-01 lk2=5.111772772e-08 wk2=1.947633683e-07 pk2=-2.568558778e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585281237e-01 ldsub=1.343555220e-11 wdsub=6.533553135e-11 pdsub=-8.616515210e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-9.109032972e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193267707e-17 nfactor=6.688221758e+00 lnfactor=-5.123670102e-07 wnfactor=-2.525315493e-06 pnfactor=3.330411325e-13 eta0=1.444049303e-02 leta0=-1.904426444e-09 weta0=-9.261004378e-09 peta0=1.221350518e-15 etab=-0.043998 u0=1.477135709e-01 lu0=-1.550569696e-08 wu0=-6.721096748e-08 pu0=8.863849602e-15 ua=-1.267244233e-09 lua=1.480064698e-17 wua=6.632216730e-17 pua=-8.746633746e-24 ub=-1.023024109e-18 lub=4.247132957e-25 wub=2.055766184e-24 pub=-2.711165001e-31 uc=2.935491635e-10 luc=-2.855819271e-17 wuc=-1.388751774e-16 puc=1.831499727e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.464148668e+05 lvsat=-2.530985185e-02 wvsat=-9.440059263e-02 pvsat=1.244964456e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000006e-02 lketa=6.282363518e-18 dwg=0.0 dwb=0.0 pclm=-2.403614773e-01 lpclm=5.536184585e-08 wpclm=2.614971561e-07 ppclm=-3.448650644e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.379922550e-24 alpha1=0.85 beta0=1.390773688e+01 lbeta0=-5.882290701e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.418817965e-01 lkt1=2.772987457e-08 wkt1=1.334169179e-07 pkt1=-1.759515655e-14 kt2=-0.028878939 at=5.372048693e+04 lat=6.915302947e-12 ute=1.528531461e-02 lute=-1.755395523e-07 wute=-8.464772511e-07 pute=1.116342663e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.108 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.109 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-8 ua=-1.245222449e-09 lua=3.748486558e-15 ub=1.918845364e-18 lub=-2.312290614e-24 wub=1.232595164e-38 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-07 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.110 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 wua=-6.617444900e-30 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917323e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 pb1=5.293955920e-35 keta=-1.740241834e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 ppclm=-1.421085472e-26 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.111 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872697e-01 leta0=-3.066156572e-7 etab=-1.378278647e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-6 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312434e-10 lb1=1.762827905e-14 keta=5.453875497e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-1 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 ub1=-1.476118686e-18 lub1=3.175805416e-24 pub1=-1.232595164e-44 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.112 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-09 peta0=6.938893904e-30 etab=7.933901887e-02 letab=-1.558362640e-07 wetab=-6.938893904e-24 petab=2.081668171e-29 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775476e-01 lags=1.437223750e-6 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 keta=6.946103312e-02 lketa=-1.257806426e-07 wketa=1.110223025e-22 pketa=-4.440892099e-28 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=-1.270549421e-26 palpha0=7.623296525e-33 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-6 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=1.654361225e-30 pua1=1.654361225e-36 ub1=9.327016030e-19 lub1=-1.525925138e-24 wub1=3.081487911e-39 pub1=-4.622231867e-45 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.113 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.308238316e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.038039511e-9 k1=6.257710814e-01 lk1=-6.813779454e-8 k2=-5.798601513e-02 lk2=2.041314719e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790972e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594373e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716768537e-9 nfactor=3.438485258e+00 lnfactor=-2.279401452e-7 eta0=-4.380244825e-01 leta0=4.193566312e-07 weta0=1.720845688e-21 peta0=-5.273559367e-28 etab=-1.600650675e-01 letab=7.204793715e-8 u0=3.089066266e-02 lu0=-2.658263485e-9 ua=-8.597024590e-10 lua=-2.657697166e-16 ub=1.904054258e-18 lub=8.862558670e-26 uc=2.781855420e-11 luc=1.116979601e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.308988651e+04 lvsat=5.742328124e-2 a0=1.033165535e+00 la0=1.588065578e-7 ags=2.238489687e+00 lags=-9.409245514e-7 a1=0.0 a2=0.42385546 b0=3.687777371e-07 lb0=-1.666436526e-13 b1=1.194667768e-08 lb1=-5.398476655e-15 keta=-1.128952678e-01 lketa=4.780085550e-08 wketa=8.881784197e-22 dwg=0.0 dwb=0.0 pclm=1.248591510e+00 lpclm=-3.600504257e-7 pdiblc1=6.447801384e-01 lpdiblc1=-2.764374541e-7 pdiblc2=8.895504641e-03 lpdiblc2=-3.998725234e-9 pdiblcb=8.513601992e-02 lpdiblcb=-8.122164671e-08 wpdiblcb=1.058181320e-22 ppdiblcb=-5.984795992e-29 drout=8.471347030e-01 ldrout=6.907687805e-8 pscbe1=1.002269402e+09 lpscbe1=-2.554584477e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094440e-06 lalpha0=-1.393643679e-12 walpha0=5.421010862e-26 alpha1=0.85 beta0=1.696331585e+01 lbeta0=4.765917258e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775674e-01 lkt1=-3.692777228e-9 kt2=-1.845629469e-02 lkt2=-8.252388786e-9 at=1.097132702e+05 lat=-4.476243271e-02 pat=2.328306437e-22 ute=-8.616208324e-01 lute=-2.027400563e-7 ua1=1.688160728e-09 lua1=-3.870320810e-16 ub1=-7.051401785e-19 lub1=3.310533463e-26 uc1=7.289584949e-11 luc1=-3.034625898e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.114 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.883840693e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.197233829e-8 k1=1.260614571e-01 lk1=1.576714902e-7 k2=8.571419420e-02 lk2=-4.452224711e-08 wk2=1.110223025e-22 pk2=8.326672685e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458427e-8 nfactor=3.214803974e+00 lnfactor=-1.268628226e-7 eta0=8.851262253e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 wetab=-4.163336342e-23 petab=-2.428612866e-29 u0=2.084392174e-02 lu0=1.881667846e-9 ua=-1.669318486e-09 lua=1.000803833e-16 wua=-1.323488980e-29 ub=2.049104468e-18 lub=2.308015275e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.493390954e+05 lvsat=3.736624816e-4 a0=1.291411731e+00 la0=4.211000822e-8 ags=-7.269793732e-01 lags=3.991145728e-7 a1=0.0 a2=0.42385546 b0=-1.068120851e-16 lb0=2.156333055e-23 b1=2.864312598e-18 lb1=-5.782502915e-25 keta=5.428652146e-02 lketa=-2.774541862e-08 wketa=-1.110223025e-22 pketa=4.163336342e-29 dwg=0.0 dwb=0.0 pclm=6.240064173e-01 lpclm=-7.781228934e-8 pdiblc1=-2.285578198e-01 lpdiblc1=1.182073759e-07 wpdiblc1=4.440892099e-22 ppdiblc1=-3.885780586e-28 pdiblc2=-6.704200072e-03 lpdiblc2=3.050484931e-09 wpdiblc2=-8.673617380e-25 ppdiblc2=6.396792818e-30 pdiblcb=-8.758737421e-02 lpdiblcb=-3.171226653e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016608e+08 lpscbe1=1.293488348e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901082e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-9 at=-3.932844299e+03 lat=6.592087176e-3 ute=-1.303201518e+00 lute=-3.198134688e-9 ua1=1.522520005e-09 lua1=-3.121821852e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=1.033975766e-31 puc1=-1.421716678e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.115 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142908321e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442105100e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220446049e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571081043e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689581891e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211731212e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135625010e-18 drout=5.033266589e-01 ldrout=1.424549367e-16 pscbe1=7.914198799e+08 lpscbe1=1.407241821e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.536504836e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610623016e-25 ub1=7.077531683e-19 lub1=2.287973959e-34 uc1=1.471862500e-10 luc1=-3.312858353e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.116 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='1.746908483e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.108198821e-08 wvth0=3.341738791e-07 pvth0=-4.407118536e-14 k1=0.90707349 k2=-2.010545839e-01 lk2=1.074764514e-08 wk2=7.631638808e-09 pk2=-1.006468158e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585275808e-01 ldsub=1.350714987e-11 wdsub=6.566741560e-11 pdsub=-8.660284435e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-9.108686028e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193267707e-17 nfactor=6.688221858e+00 lnfactor=-5.123670235e-07 wnfactor=-2.525315554e-06 pnfactor=3.330411406e-13 eta0=1.444045987e-02 leta0=-1.904422262e-09 weta0=-9.260984994e-09 peta0=1.221347962e-15 etab=-0.043998 u0=-1.478468480e-01 lu0=2.347310663e-08 wu0=1.134716189e-07 pu0=-1.496475057e-14 ua=-1.267232902e-09 lua=1.479915276e-17 wua=6.631524097e-17 pua=-8.745720294e-24 ub=-1.023024855e-18 lub=4.247133941e-25 wub=2.055766640e-24 pub=-2.711165603e-31 uc=2.946963709e-10 luc=-2.870948757e-17 wuc=-1.395764905e-16 puc=1.840748715e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.783411582e+05 lvsat=-3.144123080e-03 wvsat=8.346563073e-03 pvsat=-1.100753085e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000006e-02 lketa=6.282419029e-18 dwg=0.0 dwb=0.0 pclm=-2.403614655e-01 lpclm=5.536184429e-08 wpclm=2.614971489e-07 ppclm=-3.448650549e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.379922550e-24 alpha1=0.85 beta0=1.390773688e+01 lbeta0=-5.882290701e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.418817863e-01 lkt1=2.772987322e-08 wkt1=1.334169117e-07 pkt1=-1.759515573e-14 kt2=-0.028878939 at=5.372048693e+04 lat=6.915302947e-12 ute=2.227785078e-02 lute=-1.764617350e-07 wute=-8.507519423e-07 pute=1.121980169e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.117 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.118 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-8 ua=-1.245222449e-09 lua=3.748486558e-15 ub=1.918845364e-18 lub=-2.312290614e-24 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-07 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.119 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917323e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 keta=-1.740241833e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 wpclm=4.440892099e-22 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-08 ppdiblc2=2.775557562e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.120 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872698e-01 leta0=-3.066156572e-7 etab=-1.378278648e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-6 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312433e-10 lb1=1.762827905e-14 keta=5.453875496e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-1 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 ub1=-1.476118686e-18 lub1=3.175805416e-24 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.121 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-09 peta0=3.469446952e-30 etab=7.933901888e-02 letab=-1.558362640e-07 wetab=6.938893904e-23 petab=9.367506770e-29 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775476e-01 lags=1.437223750e-6 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 keta=6.946103312e-02 lketa=-1.257806426e-07 wketa=-5.551115123e-23 pketa=-1.665334537e-28 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=-2.752857079e-27 palpha0=1.079967008e-32 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-6 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=1.654361225e-30 pua1=-2.481541838e-36 ub1=9.327016030e-19 lub1=-1.525925138e-24 pub1=-1.540743956e-45 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.122 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='7.186223729e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.747238238e-07 wvth0=-1.129273945e-07 pvth0=1.074934412e-13 k1=6.257710822e-01 lk1=-6.813779528e-08 wk1=-4.697895406e-16 pk1=4.471836235e-22 k2=2.172676949e-02 lk2=-5.546393795e-08 wk2=-4.793305107e-08 pk2=4.562656059e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343278e-01 ldsub=4.327790950e-08 wdsub=-1.385611625e-16 pdsub=1.318953835e-22 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594364e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716769442e-09 wvoff=-5.716263018e-16 pvoff=5.441207485e-22 nfactor=3.438485268e+00 lnfactor=-2.279401540e-07 wnfactor=-5.554042559e-15 pnfactor=5.286786120e-21 eta0=-4.380244830e-01 leta0=4.193566317e-07 weta0=3.170263912e-16 peta0=-3.017719338e-22 etab=-1.600650676e-01 letab=7.204793725e-08 wetab=6.369749173e-17 petab=-6.063216595e-23 u0=-1.053975843e-02 lu0=3.677856717e-08 wu0=2.491302367e-08 pu0=-2.371423388e-14 ua=-8.597024557e-10 lua=-2.657697198e-16 wua=-1.996615475e-24 pua=1.900540102e-30 ub=1.904049007e-18 lub=8.863058489e-26 wub=3.157457102e-30 pub=-3.005523422e-36 uc=2.781855431e-11 luc=1.116979589e-17 wuc=-7.140740035e-26 puc=6.797149889e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.474474009e+05 lvsat=2.197544850e-01 wvsat=1.025478228e-01 pvsat=-9.761332408e-8 a0=1.033165529e+00 la0=1.588065632e-07 wa0=3.453642705e-15 pa0=-3.287457417e-21 ags=2.238489661e+00 lags=-9.409245272e-07 wags=1.526071713e-14 pags=-1.452638543e-20 a1=0.0 a2=0.42385546 b0=3.687777386e-07 lb0=-1.666436541e-13 wb0=-9.334353901e-22 pb0=8.885193505e-28 b1=1.194667764e-08 lb1=-5.398476615e-15 wb1=2.503135884e-23 pb1=-2.382686475e-29 keta=-1.128952687e-01 lketa=4.780085633e-08 wketa=5.265605729e-16 pketa=-5.012230631e-22 dwg=0.0 dwb=0.0 pclm=1.248591517e+00 lpclm=-3.600504321e-07 wpclm=-4.034131251e-15 ppclm=3.840014529e-21 pdiblc1=6.447801372e-01 lpdiblc1=-2.764374529e-07 wpdiblc1=7.561631321e-16 ppdiblc1=-7.197762386e-22 pdiblc2=8.895504671e-03 lpdiblc2=-3.998725263e-09 wpdiblc2=-1.822286766e-17 ppdiblc2=1.734599964e-23 pdiblcb=8.513601968e-02 lpdiblcb=-8.122164648e-08 wpdiblcb=1.464070774e-16 ppdiblcb=-1.393621199e-22 drout=8.471347039e-01 ldrout=6.907687725e-08 wdrout=-5.081908228e-16 pdrout=4.837357181e-22 pscbe1=1.002269392e+09 lpscbe1=-2.554584384e+02 wpscbe1=5.851623535e-06 ppscbe1=-5.570049286e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094428e-06 lalpha0=-1.393643668e-12 walpha0=6.868610498e-21 palpha0=-6.538077913e-27 alpha1=0.85 beta0=1.696331590e+01 lbeta0=4.765916774e-07 wbeta0=-3.058266884e-14 pbeta0=2.911104957e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775675e-01 lkt1=-3.692777150e-09 wkt1=4.907718676e-17 pkt1=-4.671640852e-23 kt2=-1.845629470e-02 lkt2=-8.252388773e-09 wkt2=7.999045870e-18 pkt2=-7.614242570e-24 at=1.097132692e+05 lat=-4.476243175e-02 wat=6.077729631e-10 pat=-5.785273388e-16 ute=-8.616208303e-01 lute=-2.027400583e-07 wute=-1.256260873e-15 pute=1.195811450e-21 ua1=1.688160724e-09 lua1=-3.870320769e-16 wua1=2.602555053e-24 pua1=-2.477323217e-30 ub1=-7.051401795e-19 lub1=3.310533553e-26 wub1=5.709966284e-34 pub1=-5.435205415e-40 uc1=7.289584960e-11 luc1=-3.034625908e-17 wuc1=-6.324064617e-26 puc1=6.019755209e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.123 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='2.127869867e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.385357636e-08 wvth0=2.258547890e-07 pvth0=-4.559579065e-14 k1=1.260614555e-01 lk1=1.576714905e-07 wk1=9.395790812e-16 pk1=-1.896833801e-22 k2=-7.371137503e-02 lk2=-1.233725376e-08 wk2=9.586610214e-08 pk2=-1.935354457e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328522e-01 ldsub=5.412372029e-08 wdsub=2.771258778e-16 pdsub=-5.594635866e-23 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994130e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458388e-08 wvoff=1.143253492e-15 pvoff=-2.308010449e-22 nfactor=3.214803955e+00 lnfactor=-1.268628188e-07 wnfactor=1.110808512e-14 pnfactor=-2.242511954e-21 eta0=8.851262263e-01 leta0=-1.785500340e-07 weta0=-6.340528103e-16 peta0=1.280033857e-22 etab=3.439973868e-02 letab=-1.582701388e-08 wetab=-1.273944422e-16 petab=2.571848810e-23 u0=1.037047639e-01 lu0=-1.484636183e-08 wu0=-4.982604734e-08 pu0=1.005893226e-14 ua=-1.669318493e-09 lua=1.000803846e-16 wua=3.993230951e-24 pua=-8.061569901e-31 ub=2.049114970e-18 lub=2.307803265e-26 wub=-6.314914204e-30 pub=1.274861193e-36 uc=2.021746669e-11 luc=1.460458297e-17 wuc=1.428150075e-25 puc=-2.883163874e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.904136703e+05 lvsat=-6.848281377e-02 wvsat=-2.050956455e-01 pvsat=4.140491401e-8 a0=1.291411743e+00 la0=4.211000591e-08 wa0=-6.907285410e-15 pa0=1.394450777e-21 ags=-7.269793224e-01 lags=3.991145626e-07 wags=-3.052143516e-14 pags=6.161697819e-21 a1=0.0 a2=0.42385546 b0=-3.211422832e-15 lb0=6.483252527e-22 wb0=1.866870744e-21 pb0=-3.768857326e-28 b1=8.611870899e-17 lb1=-1.738573109e-23 wb1=-5.006270015e-23 pb1=1.010670797e-29 keta=5.428652321e-02 lketa=-2.774541898e-08 wketa=-1.053121285e-15 pketa=2.126051557e-22 dwg=0.0 dwb=0.0 pclm=6.240064038e-01 lpclm=-7.781228663e-08 wpclm=8.068264279e-15 ppclm=-1.628829072e-21 pdiblc1=-2.285578173e-01 lpdiblc1=1.182073753e-07 wpdiblc1=-1.512324710e-15 ppdiblc1=3.053097497e-22 pdiblc2=-6.704200133e-03 lpdiblc2=3.050484943e-09 wpdiblc2=3.644574681e-17 ppdiblc2=-7.357705699e-24 pdiblcb=-8.758737372e-02 lpdiblcb=-3.171226751e-09 wpdiblcb=-2.928142173e-16 ppdiblcb=5.911360290e-23 drout=1.401075460e+00 ldrout=-1.812384256e-07 wdrout=1.016381646e-15 pdrout=-2.051878667e-22 pscbe1=1.507016803e+08 lpscbe1=1.293488309e+02 wpscbe1=-1.170324707e-05 ppscbe1=2.362663269e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901105e-06 lalpha0=-1.415246597e-12 walpha0=-1.373719389e-20 palpha0=2.773273961e-27 alpha1=0.85 beta0=2.100422365e+01 lbeta0=-1.349417754e-06 wbeta0=6.116545137e-14 pbeta0=-1.234813851e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264799e-01 lkt1=1.386230823e-08 wkt1=-9.815614987e-17 pkt1=1.981570463e-23 kt2=-4.304931438e-02 lkt2=2.860729552e-09 wkt2=-1.599831378e-17 pkt2=3.229722045e-24 at=-3.932842278e+03 lat=6.592086768e-03 wat=-1.215545519e-09 pat=2.453955531e-16 ute=-1.303201522e+00 lute=-3.198133844e-09 wute=2.512521746e-15 pute=-5.072298137e-22 ua1=1.522520013e-09 lua1=-3.121821869e-16 wua1=-5.205106796e-24 pua1=1.050812200e-30 ub1=-1.713664126e-18 lub1=4.888381450e-25 wub1=-1.141993257e-33 pub1=2.305469107e-40 uc1=-1.084804680e-10 luc1=5.161425270e-17 wuc1=1.264814733e-25 puc1=-2.553416724e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.124 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142908321e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442070405e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220668094e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571081043e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689581891e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211453656e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135402966e-18 drout=5.033266589e-01 ldrout=1.424540486e-16 pscbe1=7.914198799e+08 lpscbe1=1.407241821e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.536504836e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610623533e-25 ub1=7.077531683e-19 lub1=2.287958552e-34 uc1=1.471862500e-10 luc1=-3.312651558e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.125 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='8.609150290e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.276655848e-08 wvth0=3.874506147e-07 pvth0=-5.109737452e-14 k1=0.90707349 k2=-4.687424640e-01 lk2=4.605059045e-08 wk2=1.685982502e-07 pk2=-2.223490583e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585271307e-01 ldsub=1.356650816e-11 wdsub=6.593806449e-11 pdsub=-8.695977882e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-9.108686028e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193267707e-17 nfactor=6.688220851e+00 lnfactor=-5.123668907e-07 wnfactor=-2.525314949e-06 pnfactor=3.330410608e-13 eta0=1.444046123e-02 leta0=-1.904422441e-09 weta0=-9.260985807e-09 peta0=1.221348069e-15 etab=-0.043998 u0=1.187446795e-01 lu0=-1.168525059e-08 wu0=-4.683573157e-08 pu0=6.176743116e-15 ua=-1.267248209e-09 lua=1.480117135e-17 wua=6.632444492e-17 pua=-8.746934120e-24 ub=-1.023029542e-18 lub=4.247140122e-25 wub=2.055769459e-24 pub=-2.711169320e-31 uc=2.956530396e-10 luc=-2.883565399e-17 wuc=-1.401517565e-16 puc=1.848335380e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.734861029e+05 lvsat=-1.569193353e-02 wvsat=-4.886618534e-02 pvsat=6.444521389e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000006e-02 lketa=6.282363518e-18 dwg=0.0 dwb=0.0 pclm=-2.403614804e-01 lpclm=5.536184626e-08 wpclm=2.614971578e-07 ppclm=-3.448650667e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.379975490e-24 alpha1=0.85 beta0=1.390773688e+01 lbeta0=-5.882290701e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.418817942e-01 lkt1=2.772987426e-08 wkt1=1.334169164e-07 pkt1=-1.759515635e-14 kt2=-0.028878939 at=5.372048693e+04 lat=6.915302947e-12 ute=2.810897438e-02 lute=-1.772307494e-07 wute=-8.542583252e-07 pute=1.126604422e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.126 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.127 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-8 ua=-1.245222449e-09 lua=3.748486558e-15 ub=1.918845364e-18 lub=-2.312290614e-24 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-7 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929863e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.128 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917323e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 keta=-1.740241834e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-08 ppdiblc2=2.775557562e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 wua1=3.308722450e-30 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.129 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872698e-01 leta0=-3.066156572e-7 etab=-1.378278647e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-6 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312434e-10 lb1=1.762827905e-14 keta=5.453875497e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-1 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 pua1=6.617444900e-36 ub1=-1.476118686e-18 lub1=3.175805416e-24 pub1=3.081487911e-45 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.130 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-9 etab=7.933901888e-02 letab=-1.558362640e-07 wetab=-3.989863995e-23 petab=-6.938893904e-30 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775476e-01 lags=1.437223750e-6 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 keta=6.946103312e-02 lketa=-1.257806426e-07 wketa=-2.775557562e-23 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=-1.588186776e-27 palpha0=-1.905824131e-33 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-6 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=8.271806126e-31 pua1=4.135903063e-37 ub1=9.327016030e-19 lub1=-1.525925138e-24 pub1=-1.540743956e-45 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.131 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.243627466e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.018822352e-8 k1=6.257710813e-01 lk1=-6.813779451e-8 k2=-6.072848091e-02 lk2=2.302364826e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790973e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594374e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716768506e-9 nfactor=3.438485258e+00 lnfactor=-2.279401449e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-9.714451465e-23 peta0=-2.220446049e-28 etab=-1.600650675e-01 letab=7.204793714e-8 u0=3.231604897e-02 lu0=-4.015061633e-9 ua=-8.597024591e-10 lua=-2.657697165e-16 ub=1.904054439e-18 lub=8.862541474e-26 uc=2.781855419e-11 luc=1.116979601e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.895710940e+04 lvsat=5.183838324e-2 a0=1.033165535e+00 la0=1.588065576e-7 ags=2.238489687e+00 lags=-9.409245522e-7 a1=0.0 a2=0.42385546 b0=3.687777370e-07 lb0=-1.666436526e-13 b1=1.194667768e-08 lb1=-5.398476656e-15 keta=-1.128952678e-01 lketa=4.780085547e-8 dwg=0.0 dwb=0.0 pclm=1.248591510e+00 lpclm=-3.600504255e-7 pdiblc1=6.447801385e-01 lpdiblc1=-2.764374541e-7 pdiblc2=8.895504640e-03 lpdiblc2=-3.998725233e-9 pdiblcb=8.513601993e-02 lpdiblcb=-8.122164672e-08 wpdiblcb=-4.640385298e-23 ppdiblcb=-4.835541689e-29 drout=8.471347030e-01 ldrout=6.907687808e-8 pscbe1=1.002269402e+09 lpscbe1=-2.554584480e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094440e-06 lalpha0=-1.393643680e-12 walpha0=-1.355252716e-26 alpha1=0.85 beta0=1.696331585e+01 lbeta0=4.765917275e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775674e-01 lkt1=-3.692777231e-9 kt2=-1.845629469e-02 lkt2=-8.252388786e-9 at=1.097132703e+05 lat=-4.476243274e-2 ute=-8.616208325e-01 lute=-2.027400562e-7 ua1=1.688160728e-09 lua1=-3.870320811e-16 wua1=3.308722450e-30 ub1=-7.051401785e-19 lub1=3.310533460e-26 uc1=7.289584949e-11 luc1=-3.034625897e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.132 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.013062392e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.458107887e-8 k1=1.260614572e-01 lk1=1.576714902e-7 k2=9.119912576e-02 lk2=-4.562955058e-08 wk2=2.775557562e-23 pk2=1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458428e-8 nfactor=3.214803974e+00 lnfactor=-1.268628227e-7 eta0=8.851262252e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 wetab=1.734723476e-23 u0=1.799314912e-02 lu0=2.457184674e-9 ua=-1.669318486e-09 lua=1.000803832e-16 wua=3.308722450e-30 ub=2.049104107e-18 lub=2.308022569e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.376046496e+05 lvsat=2.742624133e-3 a0=1.291411731e+00 la0=4.211000830e-8 ags=-7.269793749e-01 lags=3.991145732e-07 wags=4.440892099e-22 pags=-3.330669074e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.428652140e-02 lketa=-2.774541861e-08 pketa=-2.081668171e-29 dwg=0.0 dwb=0.0 pclm=6.240064177e-01 lpclm=-7.781228943e-8 pdiblc1=-2.285578199e-01 lpdiblc1=1.182073759e-7 pdiblc2=-6.704200070e-03 lpdiblc2=3.050484931e-09 wpdiblc2=1.192622390e-24 ppdiblc2=-6.234162492e-31 pdiblcb=-8.758737422e-02 lpdiblcb=-3.171226649e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016602e+08 lpscbe1=1.293488349e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901081e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-9 at=-3.932844369e+03 lat=6.592087190e-03 pat=-7.275957614e-24 ute=-1.303201517e+00 lute=-3.198134717e-9 ua1=1.522520004e-09 lua1=-3.121821851e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 wub1=1.540743956e-39 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=1.292469707e-32 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.133 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142908321e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442087753e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220557072e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571063279e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689581891e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211523045e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135180921e-18 drout=5.033266589e-01 ldrout=1.424531604e-16 pscbe1=7.914198799e+08 lpscbe1=1.407337189e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.535949725e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610623275e-25 ub1=7.077531683e-19 lub1=2.287966255e-34 uc1=1.471862500e-10 luc1=-3.313065148e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.134 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='2.009340379e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.108734265e-07 wvth0=-7.305762684e-07 pvth0=9.634912886e-14 k1=0.90707349 k2=-9.090406038e-02 lk2=-3.779116058e-09 wk2=-5.104752625e-08 pk2=6.732198809e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585262889e-01 ldsub=1.367752152e-11 wdsub=6.642740346e-11 pdsub=-8.760512395e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-9.109032972e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193267707e-17 nfactor=6.688221792e+00 lnfactor=-5.123670147e-07 wnfactor=-2.525315496e-06 pnfactor=3.330411329e-13 eta0=1.444043409e-02 leta0=-1.904418861e-09 weta0=-9.260970030e-09 peta0=1.221345989e-15 etab=-0.043998 u0=-2.556520751e-01 lu0=3.769056780e-08 wu0=1.708093386e-07 pu0=-2.252650638e-14 ua=-1.267242465e-09 lua=1.480041387e-17 wua=6.632110599e-17 pua=-8.746493779e-24 ub=-1.023028196e-18 lub=4.247138347e-25 wub=2.055768676e-24 pub=-2.711168288e-31 uc=2.974364475e-10 luc=-2.907085161e-17 wuc=-1.411884907e-16 puc=1.862007934e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.808061130e+04 lvsat=1.799119811e-02 wvsat=9.960664583e-02 pvsat=-1.313622406e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000006e-02 lketa=6.282335763e-18 dwg=0.0 dwb=0.0 pclm=-2.403614720e-01 lpclm=5.536184515e-08 wpclm=2.614971529e-07 ppclm=-3.448650603e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.379975490e-24 alpha1=0.85 beta0=1.390773688e+01 lbeta0=-5.882290701e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-4.418817906e-01 lkt1=2.772987379e-08 wkt1=1.334169143e-07 pkt1=-1.759515608e-14 kt2=-0.028878939 at=5.372048693e+04 lat=6.915361155e-12 ute=3.897929900e-02 lute=-1.786643387e-07 wute=-8.605774840e-07 pute=1.134938192e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.135 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.136 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-8 ua=-1.245222449e-09 lua=3.748486558e-15 wua=6.617444900e-30 ub=1.918845364e-18 lub=-2.312290614e-24 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-7 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.137 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917322e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 keta=-1.740241834e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 wpclm=-4.440892099e-22 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 wuc1=-2.067951531e-31 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.138 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872697e-01 leta0=-3.066156572e-7 etab=-1.378278648e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-6 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312433e-10 lb1=1.762827905e-14 pb1=5.293955920e-35 keta=5.453875497e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-01 wat=9.313225746e-16 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 pua1=1.323488980e-35 ub1=-1.476118686e-18 lub1=3.175805416e-24 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.139 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-09 weta0=3.469446952e-24 peta0=3.469446952e-30 etab=7.933901888e-02 letab=-1.558362640e-07 wetab=9.367506770e-23 petab=3.989863995e-28 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775475e-01 lags=1.437223750e-06 pags=3.552713679e-27 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 keta=6.946103312e-02 lketa=-1.257806426e-07 wketa=1.665334537e-22 pketa=1.110223025e-28 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=8.470329473e-28 palpha0=5.293955920e-33 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-06 wute=1.421085472e-20 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=3.308722450e-30 pua1=4.963083675e-36 ub1=9.327016030e-19 lub1=-1.525925138e-24 wub1=1.540743956e-39 pub1=-1.540743956e-45 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.140 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.243627466e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.018822352e-8 k1=6.257710813e-01 lk1=-6.813779451e-8 k2=-6.072848091e-02 lk2=2.302364826e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790973e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594374e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716768506e-9 nfactor=3.438485258e+00 lnfactor=-2.279401449e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-3.885780586e-22 peta0=2.081668171e-28 etab=-1.600650675e-01 letab=7.204793714e-8 u0=3.231604897e-02 lu0=-4.015061633e-9 ua=-8.597024591e-10 lua=-2.657697165e-16 ub=1.904054439e-18 lub=8.862541474e-26 uc=2.781855419e-11 luc=1.116979601e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.895710940e+04 lvsat=5.183838324e-2 a0=1.033165535e+00 la0=1.588065576e-7 ags=2.238489688e+00 lags=-9.409245522e-7 a1=0.0 a2=0.42385546 b0=3.687777370e-07 lb0=-1.666436526e-13 b1=1.194667768e-08 lb1=-5.398476656e-15 keta=-1.128952678e-01 lketa=4.780085547e-8 dwg=0.0 dwb=0.0 pclm=1.248591510e+00 lpclm=-3.600504255e-7 pdiblc1=6.447801385e-01 lpdiblc1=-2.764374541e-7 pdiblc2=8.895504640e-03 lpdiblc2=-3.998725233e-9 pdiblcb=8.513601993e-02 lpdiblcb=-8.122164672e-08 wpdiblcb=3.469446952e-24 ppdiblcb=-1.994931997e-28 drout=8.471347030e-01 ldrout=6.907687808e-8 pscbe1=1.002269402e+09 lpscbe1=-2.554584480e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094440e-06 lalpha0=-1.393643680e-12 alpha1=0.85 beta0=1.696331585e+01 lbeta0=4.765917275e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775674e-01 lkt1=-3.692777231e-09 wkt1=1.776356839e-21 kt2=-1.845629469e-02 lkt2=-8.252388786e-9 at=1.097132703e+05 lat=-4.476243274e-2 ute=-8.616208325e-01 lute=-2.027400562e-7 ua1=1.688160728e-09 lua1=-3.870320811e-16 ub1=-7.051401785e-19 lub1=3.310533460e-26 uc1=7.289584949e-11 luc1=-3.034625897e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.141 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.013062392e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.458107887e-08 wvth0=3.552713679e-21 k1=1.260614572e-01 lk1=1.576714902e-7 k2=9.119912576e-02 lk2=-4.562955058e-08 pk2=-1.110223025e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458428e-8 nfactor=3.214803974e+00 lnfactor=-1.268628227e-7 eta0=8.851262252e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 petab=-2.602085214e-30 u0=1.799314912e-02 lu0=2.457184674e-9 ua=-1.669318486e-09 lua=1.000803832e-16 ub=2.049104107e-18 lub=2.308022569e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.376046496e+05 lvsat=2.742624133e-3 a0=1.291411731e+00 la0=4.211000830e-8 ags=-7.269793749e-01 lags=3.991145732e-07 wags=1.776356839e-21 pags=2.220446049e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.428652140e-02 lketa=-2.774541861e-08 wketa=-1.110223025e-22 dwg=0.0 dwb=0.0 pclm=6.240064177e-01 lpclm=-7.781228943e-8 pdiblc1=-2.285578199e-01 lpdiblc1=1.182073759e-07 ppdiblc1=-5.551115123e-29 pdiblc2=-6.704200070e-03 lpdiblc2=3.050484931e-09 wpdiblc2=-8.239936511e-24 ppdiblc2=1.734723476e-30 pdiblcb=-8.758737422e-02 lpdiblcb=-3.171226649e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016602e+08 lpscbe1=1.293488349e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901081e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-9 at=-3.932844369e+03 lat=6.592087190e-03 pat=1.455191523e-23 ute=-1.303201517e+00 lute=-3.198134717e-9 ua1=1.522520004e-09 lua1=-3.121821851e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 wub1=-6.162975822e-39 pub1=1.540743956e-45 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=-1.033975766e-31 puc1=-7.754818243e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.142 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142908321e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.796430168e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442035711e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220668094e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571081043e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689670708e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211176101e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135180921e-18 drout=5.033266589e-01 ldrout=1.424531604e-16 pscbe1=7.914198799e+08 lpscbe1=1.407241821e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.536504836e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610621982e-25 ub1=7.077531683e-19 lub1=2.287973959e-34 uc1=1.471862500e-10 luc1=-3.312858353e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.143 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-5.165351347e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.353320930e-07 wvth0=3.224989124e-06 pvth0=-4.253147906e-13 k1=0.90707349 k2=-6.220692224e-01 lk2=6.627147668e-08 wk2=2.417955132e-07 pk2=-3.188823408e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.228875002e+00 ldsub=-2.334616811e-07 wdsub=-9.759657657e-07 pdsub=1.287113411e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-9.109379917e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193178889e-17 nfactor=-1.585097167e+00 lnfactor=5.787265630e-07 wnfactor=2.035947260e-06 pnfactor=-2.685027606e-13 eta0=-9.997187851e-03 leta0=1.318439157e-09 weta0=4.212028572e-09 peta0=-5.554865401e-16 etab=-0.043998 u0=7.971402808e-01 lu0=-1.011527409e-07 wu0=-4.096182487e-07 pu0=5.402086425e-14 ua=-1.534451532e-09 lua=5.004021287e-17 wua=2.136393434e-16 pua=-2.817497024e-23 ub=3.073269759e-18 lub=-1.155100359e-25 wub=-2.026105047e-25 pub=2.672047598e-32 uc=-1.650604179e-10 luc=3.192369749e-17 wuc=1.137962061e-16 puc=-1.500755746e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.913889827e+05 lvsat=-1.103696832e-01 wvsat=-4.369996721e-01 pvsat=5.763195376e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-7.468140490e-01 lketa=9.492979659e-08 wketa=3.968493211e-07 pketa=-5.233688531e-14 dwg=0.0 dwb=0.0 pclm=1.822363870e-02 lpclm=2.125938217e-08 wpclm=1.189334925e-07 ppclm=-1.568506793e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.999997862e-08 lalpha0=2.819479502e-21 walpha0=1.179246384e-20 palpha0=-1.555201884e-27 alpha1=0.85 beta0=1.390773667e+01 lbeta0=-5.882263751e-09 wbeta0=1.126629741e-13 pbeta0=-1.485810230e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.998872425e-01 lkt1=-4.184609212e-09 wkt1=-3.935198833e-15 pkt1=5.189781938e-22 kt2=-0.028878939 at=5.372048924e+04 lat=-2.970090136e-10 wat=-1.270540990e-09 pat=1.675600652e-16 ute=-1.135968963e+00 lute=-2.371098691e-08 wute=-2.128026581e-07 pute=2.806462736e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.144 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.145 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.752573704e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.382986991e-7 k1=6.121972372e-01 lk1=-8.816639883e-7 k2=-5.601076682e-02 lk2=3.255193442e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.311152548e-7 nfactor=3.124986586e+00 lnfactor=-4.836068320e-6 eta0=0.08 etab=-0.07 u0=2.494789444e-02 lu0=3.398614506e-8 ua=-1.245222449e-09 lua=3.748486558e-15 ub=1.918845364e-18 lub=-2.312290614e-24 uc=6.326057033e-11 luc=-2.937629231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390829178e+00 la0=-5.632251912e-7 ags=3.209382116e-01 lags=4.776837126e-7 a1=0.0 a2=0.42385546 b0=6.560871865e-08 lb0=-4.269141179e-14 b1=3.134014136e-09 lb1=-1.226270809e-14 keta=-2.666112675e-03 lketa=-3.751925933e-8 dwg=0.0 dwb=0.0 pclm=-9.631270000e-03 lpclm=5.288499448e-07 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=5.528995573e-04 lpdiblc2=8.128953030e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.319501400e+07 lpscbe1=5.949551434e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832257539e-01 lkt1=-6.293314343e-8 kt2=-3.544646383e-02 lkt2=1.182853816e-7 at=1.981929862e+05 lat=-4.627437017e-1 ute=-1.016200285e+00 lute=-1.979220918e-6 ua1=1.030149760e-09 lua1=1.812633186e-15 ub1=-3.832369470e-19 lub1=-3.715699712e-24 uc1=6.920223587e-11 luc1=-7.059748407e-16 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.146 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.167677759e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.212894332e-9 k1=4.373408531e-01 lk1=5.087731700e-7 k2=1.045602503e-02 lk2=-2.030166750e-07 pk2=2.220446049e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.553724997e-9 nfactor=1.952392991e+00 lnfactor=4.488256406e-6 eta0=0.08 etab=-0.07 u0=2.778128094e-02 lu0=1.145539278e-8 ua=-9.784464677e-10 lua=1.627115701e-15 ub=1.799307847e-18 lub=-1.361742504e-24 uc=9.701328365e-12 luc=1.321337955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.408917322e+00 la0=-7.070599674e-7 ags=3.610925198e-01 lags=1.583814327e-7 a1=0.0 a2=0.42385546 b0=2.624987152e-08 lb0=2.702854569e-13 b1=-7.899974757e-10 lb1=1.894056528e-14 keta=-1.740241834e-02 lketa=7.966208966e-8 dwg=0.0 dwb=0.0 pclm=-6.899761706e-01 lpclm=5.938871634e-06 wpclm=6.661338148e-22 ppclm=6.217248938e-27 pdiblc1=0.39 pdiblc2=-1.623723774e-03 lpdiblc2=2.543720274e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.392309919e+08 lpscbe1=2.844246136e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862989458e-01 lkt1=-3.849548711e-8 kt2=-9.860889619e-03 lkt2=-8.516805990e-8 at=140000.0 ute=-1.231212620e+00 lute=-2.694684098e-7 ua1=1.514330084e-09 lua1=-2.037511139e-15 ub1=-1.026378584e-18 lub1=1.398486053e-24 uc1=-7.088796187e-11 luc1=4.080057410e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.147 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.297248088e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.299175762e-8 k1=5.592357205e-01 lk1=2.705915957e-8 k2=-3.560917656e-02 lk2=-2.097248010e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.527821500e-01 ldsub=-1.157040216e-06 wdsub=-1.776356839e-21 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.356542684e-8 nfactor=2.936087199e+00 lnfactor=6.008139587e-7 eta0=1.575872698e-01 leta0=-3.066156572e-7 etab=-1.378278647e-01 letab=2.680476500e-7 u0=3.096585297e-02 lu0=-1.129656931e-9 ua=-7.054795859e-10 lua=5.483830670e-16 ub=1.768215680e-18 lub=-1.238869957e-24 uc=3.566812735e-11 luc=2.951609590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.605932281e+00 la0=-1.485639637e-6 ags=3.277011992e-01 lags=2.903399581e-7 a1=0.0 a2=0.42385546 b0=5.038900209e-08 lb0=1.748904854e-13 b1=-4.579312434e-10 lb1=1.762827905e-14 keta=5.453875496e-04 lketa=8.734496589e-9 dwg=0.0 dwb=0.0 pclm=1.112609403e+00 lpclm=-1.184732045e-6 pdiblc1=0.39 pdiblc2=2.502894210e-03 lpdiblc2=9.129299537e-9 pdiblcb=-3.719925625e-02 lpdiblcb=4.821000899e-8 drout=0.56 pscbe1=6.245423126e+08 lpscbe1=3.424725263e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.591689679e-01 lkt1=-1.457099312e-7 kt2=-1.496516276e-02 lkt2=-6.499657985e-8 at=1.698930575e+05 lat=-1.181338060e-1 ute=-8.787696445e-01 lute=-1.662281110e-6 ua1=2.126322375e-09 lua1=-4.456031847e-15 wua1=-3.308722450e-30 ub1=-1.476118686e-18 lub1=3.175805416e-24 uc1=8.711055893e-12 luc1=9.343989506e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.148 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.816488727e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.084674858e-8 k1=5.910989287e-01 lk1=-3.513403122e-8 k2=-5.569471636e-02 lk2=1.823210342e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.567491050e-8 nfactor=3.286618135e+00 lnfactor=-8.338071560e-8 eta0=-1.433508281e-03 leta0=3.773978078e-09 peta0=-3.469446952e-30 etab=7.933901887e-02 letab=-1.558362640e-07 wetab=-2.775557562e-23 petab=3.469446952e-30 u0=3.256603176e-02 lu0=-4.253015502e-9 ua=2.554750204e-10 lua=-1.327285971e-15 pua=-1.654361225e-36 ub=3.114179744e-19 lub=1.604625805e-24 uc=6.148628680e-11 luc=-2.087787897e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.674837450e+04 lvsat=6.346786025e-3 a0=5.066918688e-01 la0=6.599468372e-7 ags=-2.598775476e-01 lags=1.437223750e-06 pags=-1.776356839e-27 a1=0.0 a2=0.42385546 b0=8.885495268e-08 lb0=9.980952730e-14 b1=1.076111291e-08 lb1=-4.269960083e-15 wb1=-2.646977960e-29 keta=6.946103312e-02 lketa=-1.257806426e-07 pketa=-8.326672685e-29 dwg=0.0 dwb=0.0 pclm=1.584889993e-01 lpclm=6.775974424e-7 pdiblc1=4.239170811e-01 lpdiblc1=-6.620210620e-8 pdiblc2=9.545914571e-03 lpdiblc2=-4.617838089e-9 pdiblcb=-2.421622557e-02 lpdiblcb=2.286867807e-8 drout=2.176050537e-01 ldrout=6.683141902e-7 pscbe1=8.629220470e+08 lpscbe1=-1.228163479e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.195826690e-06 lalpha0=1.020019183e-11 walpha0=4.870439447e-27 palpha0=4.341043855e-33 alpha1=0.85 beta0=1.042942088e+01 lbeta0=6.696082211e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.901361166e-01 lkt1=1.099223579e-7 kt2=-6.838621167e-02 lkt2=3.927495052e-8 at=1.538056803e+05 lat=-8.673316007e-2 ute=-2.354634327e+00 lute=1.218431122e-6 ua1=-1.525599643e-09 lua1=2.672085355e-15 wua1=8.271806126e-31 pua1=-2.481541838e-36 ub1=9.327016030e-19 lub1=-1.525925138e-24 wub1=7.703719778e-40 pub1=1.540743956e-45 uc1=7.140092441e-11 luc1=-2.892326820e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.149 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.243627466e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.018822352e-8 k1=6.257710813e-01 lk1=-6.813779451e-8 k2=-6.072848091e-02 lk2=2.302364826e-08 pk2=-5.551115123e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.145343276e-01 ldsub=4.327790973e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.265594374e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.716768506e-9 nfactor=3.438485258e+00 lnfactor=-2.279401449e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-3.191891196e-22 peta0=3.191891196e-28 etab=-1.600650675e-01 letab=7.204793714e-8 u0=3.231604897e-02 lu0=-4.015061633e-9 ua=-8.597024591e-10 lua=-2.657697165e-16 ub=1.904054439e-18 lub=8.862541474e-26 uc=2.781855419e-11 luc=1.116979601e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.895710940e+04 lvsat=5.183838324e-2 a0=1.033165535e+00 la0=1.588065576e-7 ags=2.238489687e+00 lags=-9.409245522e-7 a1=0.0 a2=0.42385546 b0=3.687777370e-07 lb0=-1.666436526e-13 b1=1.194667768e-08 lb1=-5.398476656e-15 keta=-1.128952678e-01 lketa=4.780085547e-8 dwg=0.0 dwb=0.0 pclm=1.248591510e+00 lpclm=-3.600504255e-7 pdiblc1=6.447801385e-01 lpdiblc1=-2.764374541e-7 pdiblc2=8.895504640e-03 lpdiblc2=-3.998725233e-9 pdiblcb=8.513601993e-02 lpdiblcb=-8.122164672e-08 wpdiblcb=5.290906602e-23 ppdiblcb=9.237402510e-29 drout=8.471347030e-01 ldrout=6.907687808e-8 pscbe1=1.002269402e+09 lpscbe1=-2.554584480e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=6.984094440e-06 lalpha0=-1.393643680e-12 alpha1=0.85 beta0=1.696331585e+01 lbeta0=4.765917275e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.707775674e-01 lkt1=-3.692777231e-9 kt2=-1.845629469e-02 lkt2=-8.252388786e-9 at=1.097132703e+05 lat=-4.476243274e-2 ute=-8.616208325e-01 lute=-2.027400562e-7 ua1=1.688160728e-09 lua1=-3.870320811e-16 ub1=-7.051401785e-19 lub1=3.310533460e-26 uc1=7.289584949e-11 luc1=-3.034625897e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.150 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.013062392e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.458107887e-8 k1=1.260614572e-01 lk1=1.576714902e-7 k2=9.119912576e-02 lk2=-4.562955058e-08 wk2=5.551115123e-23 pk2=4.857225733e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.905328527e-01 ldsub=5.412372020e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.154994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.271458428e-8 nfactor=3.214803974e+00 lnfactor=-1.268628227e-7 eta0=8.851262252e-01 leta0=-1.785500338e-7 etab=3.439973846e-02 letab=-1.582701384e-08 wetab=6.938893904e-24 petab=1.344410694e-29 u0=1.799314912e-02 lu0=2.457184674e-9 ua=-1.669318486e-09 lua=1.000803832e-16 ub=2.049104107e-18 lub=2.308022569e-26 uc=2.021746693e-11 luc=1.460458292e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.376046496e+05 lvsat=2.742624133e-3 a0=1.291411731e+00 la0=4.211000830e-8 ags=-7.269793749e-01 lags=3.991145732e-07 pags=-3.330669074e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.428652140e-02 lketa=-2.774541861e-08 wketa=2.775557562e-23 dwg=0.0 dwb=0.0 pclm=6.240064177e-01 lpclm=-7.781228943e-8 pdiblc1=-2.285578199e-01 lpdiblc1=1.182073759e-07 wpdiblc1=1.110223025e-22 ppdiblc1=-2.775557562e-29 pdiblc2=-6.704200070e-03 lpdiblc2=3.050484931e-09 wpdiblc2=-1.951563910e-24 ppdiblc2=1.111307227e-30 pdiblcb=-8.758737422e-02 lpdiblcb=-3.171226649e-9 drout=1.401075462e+00 ldrout=-1.812384259e-7 pscbe1=1.507016602e+08 lpscbe1=1.293488349e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.031901081e-06 lalpha0=-1.415246593e-12 alpha1=0.85 beta0=2.100422375e+01 lbeta0=-1.349417775e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.096264800e-01 lkt1=1.386230826e-8 kt2=-4.304931441e-02 lkt2=2.860729557e-09 wkt2=-1.110223025e-22 at=-3.932844369e+03 lat=6.592087190e-3 ute=-1.303201517e+00 lute=-3.198134717e-9 ua1=1.522520004e-09 lua1=-3.121821851e-16 ub1=-1.713664128e-18 lub1=4.888381454e-25 pub1=-3.851859889e-46 uc1=-1.084804678e-10 luc1=5.161425266e-17 wuc1=-2.584939414e-32 puc1=6.462348536e-39 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.151 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.098690578e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.630974924e-8 k1=9.070734896e-01 lk1=5.142908321e-17 k2=-1.635792203e-01 lk2=5.805356710e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-7.794653811e-18 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=5.442070405e-19 cit=0.0 voff='-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907131e-8 nfactor=2.178037929e+00 lnfactor=8.244054334e-8 eta0=2.001909455e-03 leta0=-2.640137943e-10 etab=-4.399800002e-02 letab=2.220612583e-18 u0=3.021061619e-02 lu0=-9.289795181e-12 ua=-1.208550176e-09 lua=7.060016163e-18 ub=2.099422266e-18 lub=1.292194539e-26 uc=1.218677263e-10 luc=-5.916673095e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.449528742e+05 lvsat=1.259157205e-3 a0=1.499999999e+00 la0=1.571063279e-16 ags=1.250000000e+00 lags=3.363709311e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.889316341e-01 lketa=2.135570583e-8 dwg=0.0 dwb=0.0 pclm=3.500002331e-01 lpclm=-2.249564687e-8 pdiblc1=3.569721502e-01 lpdiblc1=-2.689581891e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211592434e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135402966e-18 drout=5.033266589e-01 ldrout=1.424540486e-16 pscbe1=7.914198799e+08 lpscbe1=1.407337189e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.774280622e-09 lalpha0=3.194912098e-15 alpha1=0.85 beta0=1.518074234e+01 lbeta0=-1.737675240e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.585636645e-01 lkt1=3.553695993e-9 kt2=-2.887893901e-02 lkt2=8.535949725e-19 at=-1.837987011e+04 lat=9.508667194e-3 ute=-1.325229293e+00 lute=1.248854588e-9 ua1=-2.384733722e-11 lua1=1.610623533e-25 ub1=7.077531683e-19 lub1=2.287958552e-34 uc1=1.471862500e-10 luc1=-3.312858353e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.152 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-9.273486898e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.635035923e-08 wvth0=4.790702262e-07 pvth0=-6.318026050e-14 k1=0.90707349 k2=-2.875174805e-01 lk2=2.215045840e-08 wk2=6.069529519e-08 pk2=-8.004556225e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.238152446e+00 ldsub=-2.346851997e-07 wdsub=-9.809878504e-07 pdsub=1.293736587e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-9.109032972e-20 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.193223298e-17 nfactor=-1.585096416e+00 lnfactor=5.787264638e-07 wnfactor=2.035946853e-06 pnfactor=-2.685027069e-13 eta0=-9.997242710e-03 leta0=1.318446392e-09 weta0=4.212058269e-09 peta0=-5.554904565e-16 etab=-0.043998 u0=4.727431475e-02 lu0=-2.259667426e-09 wu0=-3.699304184e-09 pu0=4.878679351e-16 ua=-1.534448332e-09 lua=5.003979081e-17 wua=2.136376110e-16 pua=-2.817474177e-23 ub=3.073243389e-18 lub=-1.155065582e-25 wub=-2.025962301e-25 pub=2.671859343e-32 uc=-1.661421677e-10 luc=3.206635973e-17 wuc=1.143817810e-16 puc=-1.508478367e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.670452138e+05 lvsat=-1.484250264e-02 wvsat=-4.489645444e-02 pvsat=5.920989308e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-7.468145630e-01 lketa=9.492986439e-08 wketa=3.968495993e-07 pketa=-5.233692201e-14 dwg=0.0 dwb=0.0 pclm=1.822366269e-02 lpclm=2.125937901e-08 wpclm=1.189334796e-07 ppclm=-1.568506622e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-1.998733058e-24 walpha0=2.113544139e-22 palpha0=-2.787363083e-29 alpha1=0.85 beta0=1.390773688e+01 lbeta0=-5.882291190e-09 wbeta0=3.831246431e-17 pbeta0=-5.059064279e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.998872496e-01 lkt1=-4.184608273e-09 wkt1=-7.863398821e-17 pkt1=1.037037123e-23 kt2=-0.028878939 at=5.372048694e+04 lat=6.448710337e-12 wat=-2.496084198e-11 pat=3.291876055e-18 ute=-1.133946109e+00 lute=-2.397776296e-08 wute=-2.138976737e-07 pute=2.820903910e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.153 nmos lmin=2.0e-05 lmax=0.0001 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.154 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.490906710e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.603735711e-07 wvth0=1.364127605e-08 pvth0=-2.721691164e-13 k1=8.459775980e-01 lk1=-5.546021926e-06 wk1=-1.218748452e-07 pk1=2.431632409e-12 k2=-1.555260221e-01 lk2=2.311035875e-06 wk2=5.187949190e-08 pk2=-1.035093449e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.013920080e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.373853003e-07 wvoff=-1.638297997e-10 pvoff=3.268712669e-15 nfactor=3.855575864e+00 lnfactor=-1.941269866e-05 wnfactor=-3.808722637e-07 pnfactor=7.599118081e-12 eta0=0.08 etab=-0.07 u0=2.216136417e-02 lu0=8.958266540e-08 wu0=1.452679533e-09 pu0=-2.898368917e-14 ua=-1.666460410e-09 lua=1.215297622e-14 wua=2.196006162e-16 pua=-4.381445361e-21 ub=2.233762623e-18 lub=-8.595482281e-24 wub=-1.641732951e-25 pub=3.275566046e-30 uc=6.321310771e-11 luc=-2.928159546e-16 wuc=2.474330664e-20 puc=-4.936755097e-25 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.022295913e+00 la0=6.789706651e-06 wa0=1.921244986e-07 pa0=-3.833245134e-12 ags=3.185092424e-01 lags=5.261462180e-07 wags=1.266275105e-09 pags=-2.526457020e-14 a1=0.0 a2=0.42385546 b0=1.200539247e-07 lb0=-1.128975683e-12 wb0=-2.838348370e-14 pb0=5.663038891e-19 b1=4.708097883e-09 lb1=-4.366863971e-14 wb1=-8.206044874e-16 pb1=1.637260308e-20 keta=-5.571941629e-03 lketa=2.045749416e-08 wketa=1.514872562e-09 pketa=-3.022455709e-14 dwg=0.0 dwb=0.0 pclm=6.479011413e-02 lpclm=-9.559966552e-07 wpclm=-3.879750482e-08 ppclm=7.740831992e-13 pdiblc1=0.39 pdiblc2=3.520759640e-03 lpdiblc2=-5.108543816e-08 wpdiblc2=-1.547210754e-09 ppdiblc2=3.086976484e-14 pdiblcb=-0.025 drout=0.56 pscbe1=-1.067736711e+08 lpscbe1=6.619508806e+03 wpscbe1=1.750529270e+01 ppscbe1=-3.492635168e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.029925381e-01 lkt1=3.314513827e-07 wkt1=1.030485947e-08 pkt1=-2.056013299e-13 kt2=-6.483309138e-02 lkt2=7.046038775e-07 wkt2=1.531989545e-08 pkt2=-3.056607309e-13 at=2.400717663e+05 lat=-1.298304138e+00 wat=-2.183232939e-02 pat=4.355960380e-7 ute=-5.625135003e-01 lute=-1.103112565e-05 wute=-2.365169017e-07 pute=4.718957078e-12 ua1=1.673407822e-09 lua1=-1.102157512e-14 wua1=-3.353445794e-16 pua1=6.690755143e-21 ub1=-9.468974077e-19 lub1=7.530386725e-24 wub1=2.938485987e-25 pub1=-5.862832274e-30 uc1=1.790432795e-10 luc1=-2.897510272e-15 wuc1=-5.726255254e-17 puc1=1.142495634e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.155 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.179237923e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=3.130207820e-07 wvth0=-6.026567759e-10 pvth0=-1.589030576e-13 k1=-2.781159300e-01 lk1=3.392636040e-06 wk1=3.729833611e-07 pk1=-1.503421159e-12 k2=3.123990654e-01 lk2=-1.409848737e-06 wk2=-1.574095497e-07 pk2=6.291481045e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.451672935e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.715755081e-07 wvoff=-1.745528365e-08 pvoff=1.407682960e-13 nfactor=-2.910718754e-01 lnfactor=1.356095072e-05 wnfactor=1.169567591e-06 pnfactor=-4.729795143e-12 eta0=0.08 etab=-0.07 u0=3.250448028e-02 lu0=7.335436892e-09 wu0=-2.462307728e-09 pu0=2.147823643e-15 ua=1.007938084e-10 lua=-1.900019016e-15 wua=-5.626316992e-16 pua=1.838772925e-21 ub=8.062373536e-19 lub=2.756028785e-24 wub=5.177094959e-25 pub=-2.146684764e-30 uc=-8.646487960e-11 luc=8.974055888e-16 wuc=5.013355987e-17 puc=-3.989530219e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.264764956e+00 la0=-3.090259324e-06 wa0=-4.461721998e-07 pa0=1.242414255e-12 ags=1.701178370e-01 lags=1.706137015e-06 wags=9.955930356e-08 pags=-8.068790356e-13 a1=0.0 a2=0.42385546 b0=-2.767762927e-07 lb0=2.026570983e-12 wb0=1.579742060e-13 pb0=-9.155902829e-19 b1=1.287408912e-08 lb1=-1.086036303e-13 wb1=-7.123388953e-15 pb1=6.649159512e-20 keta=-9.931611010e-03 lketa=5.512506628e-08 wketa=-3.894696216e-09 pketa=1.279169010e-14 dwg=0.0 dwb=0.0 pclm=-2.153176552e+00 lpclm=1.668101033e-05 wpclm=7.627985490e-07 ppclm=-5.600113231e-12 pdiblc1=0.39 pdiblc2=-4.145556882e-03 lpdiblc2=9.876198533e-09 wpdiblc2=1.314687080e-09 ppdiblc2=8.112293836e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.109587882e+09 lpscbe1=-3.052853519e+03 wpscbe1=-2.452073947e+02 ppscbe1=1.739796511e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.009252328e-01 lkt1=3.150124174e-07 wkt1=7.625005222e-09 pkt1=-1.842914478e-13 kt2=2.715659367e-02 lkt2=-2.688715133e-08 wkt2=-1.929802843e-08 pkt2=-3.038311981e-14 at=1.436365975e+04 lat=4.964998659e-01 wat=6.549698817e-02 pat=-2.588363031e-7 ute=-3.011856604e+00 lute=8.445759237e-06 wute=9.282888826e-07 pute=-4.543439907e-12 ua1=-2.164666612e-09 lua1=1.949833605e-14 wua1=1.917941916e-15 pua1=-1.122711093e-20 ub1=1.746654036e-18 lub1=-1.388841382e-23 wub1=-1.445642911e-24 pub1=7.969397215e-30 uc1=-3.198216898e-10 luc1=1.069404599e-15 wuc1=1.297746289e-16 puc1=-3.448017754e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.156 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.281322442e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.225099051e-07 wvth0=-5.130196107e-08 pvth0=4.145455971e-14 k1=7.140556678e-01 lk1=-5.283080456e-07 wk1=-8.071104457e-08 pk1=2.895251421e-13 k2=-9.638710442e-02 lk2=2.056255599e-07 wk2=3.168487091e-08 pk2=-1.181305434e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.086337760e+00 ldsub=-6.031905193e-06 wdsub=-6.430796777e-07 pdsub=2.541374360e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.441888683e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.594297841e-07 wvoff=5.587578944e-08 pvoff=-1.490273784e-13 nfactor=3.880766189e+00 lnfactor=-2.925656866e-06 wnfactor=-4.924819408e-07 pnfactor=1.838426823e-12 eta0=4.844795064e-01 leta0=-1.598454876e-06 weta0=-1.704161146e-07 peta0=6.734642054e-13 etab=-4.236015811e-01 letab=1.397391370e-06 wetab=1.489801253e-07 petab=-5.887517267e-13 u0=3.669216835e-02 lu0=-9.213808019e-09 wu0=-2.985254186e-09 pu0=4.214445814e-15 ua=-1.593280350e-09 lua=4.794760465e-15 wua=4.628300702e-16 pua=-2.213729958e-21 ub=3.521107115e-18 lub=-7.972813442e-24 wub=-9.138208688e-25 pub=3.510552886e-30 uc=2.063485884e-10 luc=-2.597583919e-16 wuc=-8.897947931e-17 puc=1.508051545e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.596059383e+05 lvsat=-1.104969395e+00 wvsat=-1.457647270e-01 pvsat=5.760448549e-7 a0=4.799522055e+00 la0=-1.310731774e-05 wa0=-1.664888608e-06 pa0=6.058636474e-12 ags=-1.313286725e-01 lags=2.897417748e-06 wags=2.393023707e-07 pags=-1.359127008e-12 a1=0.0 a2=0.42385546 b0=5.752437132e-08 lb0=7.054545400e-13 wb0=-3.719824961e-15 pb0=-2.765947141e-19 b1=-4.424871597e-08 lb1=1.171388978e-13 wb1=2.282909948e-14 pb1=-5.187707481e-20 keta=5.610142409e-02 lketa=-2.058296305e-07 wketa=-2.896258408e-08 pketa=1.118569999e-13 dwg=0.0 dwb=0.0 pclm=8.904007843e+00 lpclm=-2.701566659e-05 wpclm=-4.061827418e-06 ppclm=1.346623446e-11 pdiblc1=0.39 pdiblc2=1.537764194e-02 lpdiblc2=-6.727715993e-08 wpdiblc2=-6.711889234e-09 ppdiblc2=3.983236826e-14 pdiblcb=-8.859740667e-02 lpdiblcb=2.513293831e-07 wpdiblcb=2.679498657e-08 ppdiblcb=-1.058905983e-13 drout=0.56 pscbe1=-1.146995250e+08 lpscbe1=1.785384624e+03 wpscbe1=3.853830333e+02 ppscbe1=-7.522218203e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-6.275471608e-02 lkt1=-6.262091225e-07 wkt1=-1.023950706e-07 pkt1=2.504947994e-13 kt2=1.606047841e-01 lkt2=-5.542585197e-07 wkt2=-9.152847585e-08 pkt2=2.550630130e-13 at=2.958390853e+05 lat=-6.158575202e-01 wat=-6.565843510e-02 pat=2.594743221e-7 ute=2.203824086e+00 lute=-1.216599018e-05 wute=-1.607023929e-06 pute=5.475814621e-12 ua1=1.240858312e-08 lua1=-3.809341267e-14 wua1=-5.360368735e-15 pua1=1.753590665e-20 ub1=-7.928595002e-18 lub1=2.434701902e-23 wub1=3.363817858e-24 pub1=-1.103701942e-29 uc1=-1.991689359e-10 luc1=5.925992733e-16 wuc1=1.083724131e-16 puc1=-2.602227654e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.157 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.706409780e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.848943050e-07 wvth0=5.738657666e-09 pvth0=-6.988194022e-14 k1=4.639892783e-01 lk1=-4.020821110e-08 wk1=6.626505721e-08 pk1=2.645281601e-15 k2=-1.965783151e-02 lk2=5.585914999e-08 wk2=-1.878682088e-08 pk2=-1.961580717e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-2.207111220e+00 ldsub=2.348396295e-06 wdsub=1.286159355e-06 pdsub=-1.224270653e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='7.154520925e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.568455630e-07 wvoff=-7.153405026e-08 pvoff=9.966146688e-14 nfactor=3.706128668e+00 lnfactor=-2.584785206e-06 wnfactor=-2.187000700e-07 pnfactor=1.304037192e-12 eta0=-6.552179816e-01 leta0=6.260989963e-07 weta0=3.408322292e-07 peta0=-3.244317232e-13 etab=9.880177684e-01 letab=-1.357921618e-06 wetab=-4.737142231e-07 petab=6.266735407e-13 u0=2.689597896e-02 lu0=9.907187920e-09 wu0=2.955923264e-09 pu0=-7.382025568e-15 ua=2.402332641e-09 lua=-3.004200617e-15 wua=-1.119204109e-15 pua=8.742124970e-22 ub=-3.316125579e-18 lub=5.372651145e-24 wub=1.891118260e-24 pub=-1.964354506e-30 uc=1.173430744e-10 luc=-8.603022019e-17 wuc=-2.911937222e-17 puc=3.396534883e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.111568452e+05 lvsat=-1.860964624e-01 wvsat=9.795912495e-02 pvsat=1.003248991e-7 a0=-3.678333816e+00 la0=3.440448051e-06 wa0=2.181745960e-06 pa0=-1.449536454e-12 ags=-2.750675914e+00 lags=8.010071861e-06 wags=1.298507986e-06 pags=-3.426570323e-12 a1=0.0 a2=0.42385546 b0=-6.464351611e-07 lb0=2.079499776e-12 wb0=3.833229127e-13 pb0=-1.032056080e-18 b1=3.726031130e-08 lb1=-4.195702383e-14 wb1=-1.381461510e-14 pb1=1.964709545e-20 keta=2.860668266e-01 lketa=-6.546947304e-07 wketa=-1.129213655e-07 pketa=2.757345501e-13 dwg=0.0 dwb=0.0 pclm=-9.802592466e+00 lpclm=9.497391129e-06 wpclm=5.192930912e-06 ppclm=-4.597952484e-12 pdiblc1=1.366529826e+00 lpdiblc1=-1.906070014e-06 wpdiblc1=-4.914047615e-07 ppdiblc1=9.591636174e-13 pdiblc2=-3.714385982e-02 lpdiblc2=3.523856143e-08 wpdiblc2=2.434040656e-08 ppdiblc2=-2.077801791e-14 pdiblcb=-2.091401144e-02 lpdiblcb=1.192194499e-07 wpdiblcb=-1.721516871e-09 ppdiblcb=-5.022977707e-14 drout=-8.470974543e-01 ldrout=2.746486786e-06 wdrout=5.550528409e-07 pdrout=-1.083397094e-12 pscbe1=1.128026474e+09 lpscbe1=-6.402686414e+02 wpscbe1=-1.382047699e+02 ppscbe1=2.697592645e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.721338422e-05 lalpha0=5.317584403e-11 walpha0=1.147823713e-11 palpha0=-2.240415296e-17 alpha1=0.85 beta0=-4.024363701e+00 lbeta0=3.490814970e-05 wbeta0=7.535075883e-06 pbeta0=-1.470757145e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-5.727589350e-01 lkt1=3.692584223e-07 wkt1=9.520529294e-08 pkt1=-1.351975958e-13 kt2=-2.122811782e-01 lkt2=1.735705054e-07 wkt2=7.501561177e-08 pkt2=-7.001122729e-14 at=1.718672079e+05 lat=-3.738791682e-01 wat=-9.415871704e-03 pat=1.496955313e-7 ute=-5.415833772e+00 lute=2.706675218e-06 wute=1.595870617e-06 pute=-7.758543886e-13 ua1=-1.143250815e-08 lua1=8.441560401e-15 wua1=5.164689358e-15 pua1=-3.007754270e-21 ub1=6.732271364e-18 lub1=-4.269247481e-24 wub1=-3.023443307e-24 pub1=1.430154290e-30 uc1=1.910574971e-10 luc1=-1.690762871e-16 wuc1=-6.237960380e-17 puc1=7.306485212e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.158 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.811588157e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.549362488e-08 wvth0=-8.174124034e-08 pvth0=1.338851257e-14 k1=7.563678524e-01 lk1=-3.185178206e-07 wk1=-6.808296987e-08 pk1=1.305286160e-13 k2=-6.280301337e-02 lk2=9.692822884e-08 wk2=1.081499412e-09 pk2=-3.852808376e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.951761930e-01 ldsub=6.170455024e-08 wdsub=1.009182144e-08 pdsub=-9.606213081e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.076008340e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.868251810e-09 wvoff=4.224866296e-08 pvoff=-8.646135961e-15 nfactor=1.101542506e+00 lnfactor=-1.055291262e-07 wnfactor=1.218299669e-06 pnfactor=-6.381555709e-14 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-2.775557562e-23 peta0=-4.683753385e-29 etab=-8.331377799e-01 letab=3.756017469e-07 wetab=3.508876126e-07 petab=-1.582492792e-13 u0=5.984836800e-02 lu0=-2.145956511e-08 wu0=-1.435320362e-08 pu0=9.094203443e-15 ua=9.451187017e-10 lua=-1.617106355e-15 wua=-9.408929772e-16 pua=7.044815190e-22 ub=1.426680081e-18 lub=8.580645503e-25 wub=2.488657547e-25 pub=-4.011255490e-31 uc=-1.794271043e-10 luc=1.964596743e-16 wuc=1.080417212e-16 puc=-9.659568993e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-7.194896744e+05 lvsat=3.929639994e-01 wvsat=3.901817742e-01 pvsat=-1.778362885e-7 a0=-9.337107707e-01 la0=8.278935221e-07 wa0=1.025375889e-06 pa0=-3.488097545e-13 ags=1.012170807e+01 lags=-4.242905873e-06 wags=-4.109695171e-06 pags=1.721395506e-12 a1=0.0 a2=0.42385546 b0=2.928340857e-06 lb0=-1.323261595e-12 wb0=-1.334356565e-12 pb0=6.029703789e-19 b1=-1.297928289e-08 lb1=5.865091333e-15 wb1=1.299445162e-14 pb1=-5.871945791e-21 keta=-7.379365300e-01 lketa=3.200346087e-07 wketa=3.258477609e-07 pketa=-1.419214447e-13 dwg=0.0 dwb=0.0 pclm=5.695165307e-01 lpclm=-3.756223553e-07 wpclm=3.540167263e-07 ppclm=8.117989621e-15 pdiblc1=5.364444156e-01 lpdiblc1=-1.115927483e-06 wpdiblc1=5.647779571e-08 ppdiblc1=4.376446209e-13 pdiblc2=4.590637652e-03 lpdiblc2=-4.487713755e-09 wpdiblc2=2.244221868e-09 ppdiblc2=2.549204742e-16 pdiblcb=5.491633018e-01 lpdiblcb=-4.234263131e-07 wpdiblcb=-2.419076307e-07 ppdiblcb=1.783988211e-13 drout=2.976540100e+00 ldrout=-8.931611524e-07 wdrout=-1.110105880e-06 pdrout=5.016358545e-13 pscbe1=1.854474894e+09 lpscbe1=-1.331761090e+03 wpscbe1=-4.442734713e+02 ppscbe1=5.611002461e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.845364065e-05 lalpha0=-9.331349271e-12 walpha0=-1.640576677e-11 palpha0=4.138100554e-18 alpha1=0.85 beta0=3.666375002e+01 lbeta0=-3.822092671e-06 wbeta0=-1.027026974e-05 pbeta0=2.240998748e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.020959911e-01 lkt1=1.643140867e-08 wkt1=-3.580521670e-08 pkt1=-1.049118084e-14 kt2=-7.392936336e-02 lkt2=4.187604154e-08 wkt2=2.891933110e-08 pkt2=-2.613305355e-14 at=-4.707664425e+05 lat=2.378315935e-01 wat=3.026168448e-01 pat=-1.473224830e-7 ute=-4.376328549e+00 lute=1.717189947e-06 wute=1.832294456e-06 pute=-1.000901749e-12 ua1=-7.358206390e-09 lua1=4.563309965e-15 wua1=4.716070199e-15 pua1=-2.580722216e-21 ub1=7.457050586e-18 lub1=-4.959151052e-24 wub1=-4.255129614e-24 pub1=2.602573084e-30 uc1=4.033700770e-10 luc1=-3.711725979e-16 wuc1=-1.722834852e-16 puc1=1.776802687e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.159 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='7.819915037e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.105800074e-08 wvth0=-9.419520343e-08 pvth0=1.901622186e-14 k1=-6.394018493e-01 lk1=3.122039879e-07 wk1=3.990528618e-07 pk1=-8.056119080e-14 k2=3.830676809e-01 lk2=-1.045522664e-07 wk2=-1.521574989e-07 pk2=3.071770803e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.292491219e-01 ldsub=4.630764106e-08 wdsub=-2.018364287e-08 pdsub=4.074694007e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590353e-03 lcdscd=-1.221701112e-9 cit=0.0 voff='-1.956435991e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.465004556e-09 wvoff=4.178092842e-08 pvoff=-8.434775610e-15 nfactor=-5.196320614e-01 lnfactor=6.270488586e-07 wnfactor=1.946843663e-06 pnfactor=-3.930307455e-13 eta0=8.851262252e-01 leta0=-1.785500338e-7 etab=3.201989587e-02 letab=-1.534656884e-08 wetab=1.240664295e-09 petab=-2.504665486e-16 u0=-2.019537367e-03 lu0=6.497365835e-09 wu0=1.043305374e-08 pu0=-2.106235323e-15 ua=-3.812407475e-09 lua=5.327293315e-16 wua=1.117239438e-15 pua=-2.255494150e-22 ub=4.263995041e-18 lub=-4.240641710e-25 wub=-1.154671372e-24 pub=2.331062112e-31 uc=3.867754784e-10 luc=-5.939651500e-17 wuc=-1.910947557e-16 puc=3.857840037e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.492715899e+05 lvsat=3.872905620e-04 wvsat=-6.082232641e-03 pvsat=1.227887208e-9 a0=4.125834615e-01 la0=2.195287381e-07 wa0=4.581525110e-07 pa0=-9.249228707e-14 ags=3.142017554e-01 lags=1.889198854e-07 wags=-5.427906292e-07 pags=1.095791150e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.344445194e-02 lketa=-1.950018079e-08 wketa=2.129186933e-08 pketa=-4.298423872e-15 dwg=0.0 dwb=0.0 pclm=-6.657256243e-01 lpclm=1.825601049e-07 wpclm=6.723656876e-07 ppclm=-1.357378574e-13 pdiblc1=-3.782337355e+00 lpdiblc1=8.356479422e-07 wpdiblc1=1.852663455e-06 ppdiblc1=-3.740175509e-13 pdiblc2=-1.644130456e-02 lpdiblc2=5.016221321e-09 wpdiblc2=5.076166784e-09 ppdiblc2=-1.024781627e-15 pdiblcb=-6.176655912e-01 lpdiblcb=1.038414939e-07 wpdiblcb=2.763414362e-07 ppdiblcb=-5.578808548e-14 drout=1.401074700e+00 ldrout=-1.812382722e-07 wdrout=3.970125744e-13 pdrout=-8.014929553e-20 pscbe1=-2.614127030e+09 lpscbe1=6.875152157e+02 wpscbe1=1.441366022e+03 ppscbe1=-2.909844140e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.216303876e-05 lalpha0=-6.488745799e-12 walpha0=-1.310141496e-11 palpha0=2.644926753e-18 alpha1=0.85 beta0=3.941849373e+01 lbeta0=-5.066909012e-06 wbeta0=-9.599764052e-06 pbeta0=1.938009966e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.049861390e-01 lkt1=-2.745068843e-08 wkt1=-1.066835119e-07 pkt1=2.153737406e-14 kt2=5.719550391e-02 lkt2=-1.737679461e-08 wkt2=-5.225982918e-08 pkt2=1.055026657e-14 at=7.721224839e+04 lat=-9.789565281e-03 wat=-4.230272205e-02 pat=8.540115829e-9 ute=2.359994270e-02 lute=-2.710541403e-07 wute=-6.916907908e-07 pute=1.396392285e-13 ua1=4.972362508e-09 lua1=-1.008639840e-15 wua1=-1.798478793e-15 pua1=3.630786973e-22 ub1=-6.929333973e-18 lub1=1.541782789e-24 wub1=2.719043435e-24 pub1=-5.489232077e-31 uc1=-8.744457260e-10 luc1=2.062480850e-16 wuc1=3.993145404e-16 puc1=-8.061401872e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.160 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='3.652038560e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.308350636e-08 wvth0=1.275493523e-07 pvth0=-2.574979079e-14 k1=9.070734896e-01 lk1=5.142886117e-17 k2=-2.559449716e-01 lk2=2.445224694e-08 wk2=4.815229817e-08 pk2=-9.721034107e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.769155277e+00 ldsub=-2.645701535e-07 wdsub=-6.832056585e-07 pdsub=1.379262415e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999994e-03 lcdscd=8.701208157e-19 wcdscd=8.416132374e-19 pcdscd=-1.699055393e-25 cit=0.0 voff='-1.237493846e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.104907135e-08 wvoff=-1.102522518e-16 pvoff=2.225786222e-23 nfactor=-5.352926522e+00 lnfactor=1.602799178e-06 wnfactor=3.926057449e-06 pnfactor=-7.925964039e-13 eta0=2.001908064e-03 leta0=-2.640134732e-10 weta0=8.292438567e-16 peta0=-1.674085790e-22 etab=-4.399800002e-02 letab=2.220570949e-18 u0=-6.625188931e-03 lu0=7.427159378e-09 wu0=1.920331560e-08 pu0=-3.876784556e-15 ua=-1.256820177e-09 lua=1.680481206e-17 wua=2.516421301e-17 pua=-5.080176487e-24 ub=2.699802203e-18 lub=-1.082833566e-25 wub=-3.129912694e-25 pub=6.318699046e-32 uc=2.366081437e-10 luc=-2.908058330e-17 wuc=-5.981670388e-17 puc=1.207585600e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.301128123e+05 lvsat=4.255083741e-03 wvsat=7.736450749e-03 pvsat=-1.561842414e-9 a0=1.499999999e+00 la0=1.571063279e-16 ags=1.250000000e+00 lags=3.363798129e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.173646676e-01 lketa=8.766009508e-08 wketa=1.712193659e-07 pketa=-3.456593681e-14 dwg=0.0 dwb=0.0 pclm=3.636937568e-01 lpclm=-2.526010913e-08 wpclm=-7.138735169e-09 ppclm=1.441174995e-15 pdiblc1=3.569721502e-01 lpdiblc1=-2.689626299e-17 pdiblc2=8.406112095e-03 lpdiblc2=7.211488351e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.135264188e-18 drout=5.033266589e-01 ldrout=1.424536045e-16 pscbe1=7.914198799e+08 lpscbe1=1.407337189e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.772300406e-07 lalpha0=-3.141874819e-14 walpha0=-8.938365973e-14 palpha0=1.804486261e-20 alpha1=0.85 beta0=1.944226051e+01 lbeta0=-1.034087074e-06 wbeta0=-2.221623175e-06 pbeta0=4.485035083e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.739733244e-01 lkt1=-1.352348645e-08 wkt1=-4.409880527e-08 pkt1=8.902710907e-15 kt2=-2.887893901e-02 lkt2=8.536088503e-19 at=-9.775753668e+04 lat=2.553350990e-02 wat=4.138132389e-02 pat=-8.354103048e-9 ute=-1.033781996e+00 lute=-5.758881717e-08 wute=-1.519378877e-07 pute=3.067337272e-14 ua1=-2.384733722e-11 lua1=1.610623275e-25 ub1=7.077531683e-19 lub1=2.287968181e-34 uc1=1.471862500e-10 luc1=-3.312858353e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.161 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='1.272009734e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.650695965e-08 wvth0=-2.324011598e-07 pvth0=2.172084269e-14 k1=0.90707349 k2=2.156852212e-02 lk2=-1.214651012e-08 wk2=-1.004380379e-07 pk2=9.875208001e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-7.698091194e-01 ldsub=7.027101011e-08 wdsub=5.871286889e-07 pdsub=-2.960672252e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000005e-03 lcdscd=-4.748623370e-19 wcdscd=-1.963762486e-18 pcdscd=2.000704290e-25 cit=0.0 voff='-2.075300006e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.220768345e-17 wvoff=2.572555502e-16 pvoff=-2.620942352e-23 nfactor=1.598715371e+01 lnfactor=-1.211551944e-06 wnfactor=-7.124853728e-06 pnfactor=6.648088131e-13 eta0=-9.997241958e-03 leta0=1.318446536e-09 weta0=4.212058397e-09 peta0=-5.554905315e-16 etab=-0.043998 u0=6.352376718e-02 lu0=-1.824155103e-09 wu0=-1.217050122e-08 pu0=2.608257799e-16 ua=-1.421817344e-09 lua=3.856480353e-17 wua=1.549205992e-16 pua=-2.219257845e-23 ub=1.672391278e-18 lub=2.721262354e-26 wub=5.276987942e-25 pub=-4.768405582e-32 uc=-4.396916632e-10 luc=6.011051154e-17 wuc=2.569891512e-16 puc=-2.970481697e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.747358051e+05 lvsat=-1.481794118e-02 wvsat=-4.890572889e-02 pvsat=5.908184879e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.952945678e-02 lketa=1.685396106e-08 wketa=-2.662397749e-09 pketa=-1.163423594e-14 dwg=0.0 dwb=0.0 pclm=-1.372788984e-02 lpclm=2.451463505e-08 wpclm=1.355905268e-07 ppclm=-1.738210281e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.700634379e-07 lalpha0=4.075886305e-14 walpha0=2.085618718e-13 palpha0=-2.124849203e-20 alpha1=0.85 beta0=3.964194500e+00 lbeta0=1.007175750e-06 wbeta0=5.183787401e-06 pbeta0=-5.281294439e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.972647105e-01 lkt1=1.592440484e-08 wkt1=1.028972126e-07 pkt1=-1.048327093e-14 kt2=-0.028878939 at=2.389350420e+05 lat=-1.886984407e-02 wat=-9.655642231e-02 pat=9.837264859e-9 ute=-1.803102747e+00 lute=4.386997276e-08 wute=1.349484029e-07 pute=-7.161478179e-15 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.162 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.163 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.814679883e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.143851906e-7 k1=5.567098995e-01 lk1=2.254127697e-7 k2=-3.239100444e-02 lk2=-1.457393440e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017808550e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.296270710e-7 nfactor=2.951582568e+00 lnfactor=-1.376331981e-6 eta0=0.08 etab=-0.07 u0=2.560927226e-02 lu0=2.079041345e-8 ua=-1.145242396e-09 lua=1.753696429e-15 ub=1.844100334e-18 lub=-8.209866543e-25 uc=6.327183549e-11 luc=-2.939876843e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.478299869e+00 la0=-2.308430009e-6 ags=3.215147230e-01 lags=4.661812263e-7 a1=0.0 a2=0.42385546 b0=5.268624936e-08 lb0=2.151361575e-13 b1=2.760408260e-09 lb1=-4.808568123e-15 wb1=-3.308722450e-30 keta=-1.976419529e-03 lketa=-5.127993490e-8 dwg=0.0 dwb=0.0 pclm=-2.729504833e-02 lpclm=8.812755480e-07 ppclm=2.220446049e-28 pdiblc1=0.39 pdiblc2=-1.515165620e-04 lpdiblc2=2.218337962e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.522518163e+07 lpscbe1=5.790538287e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.785341441e-01 lkt1=-1.565395837e-7 kt2=-2.847160196e-02 lkt2=-2.087623258e-8 at=1.882531350e+05 lat=-2.644249724e-1 ute=-1.123882006e+00 lute=1.692319823e-7 ua1=8.774736444e-10 lua1=4.858808868e-15 ub1=-2.494531757e-19 lub1=-6.384937596e-24 uc1=4.313166665e-11 luc1=-1.858179462e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.164 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.164933975e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-6.413269591e-8 k1=6.071532016e-01 lk1=-1.757063659e-7 k2=-6.120959896e-02 lk2=8.342269022e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.259465233e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.253544744e-8 nfactor=2.484875242e+00 lnfactor=2.334869137e-6 eta0=0.08 etab=-0.07 u0=2.666023828e-02 lu0=1.243325671e-8 ua=-1.234602158e-09 lua=2.464274623e-15 ub=2.035011298e-18 lub=-2.339087928e-24 uc=3.252620055e-11 luc=-4.950205394e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.205783464e+00 la0=-1.414119935e-7 ags=4.064200087e-01 lags=-2.089755015e-7 a1=0.0 a2=0.42385546 b0=9.817257298e-08 lb0=-1.465656750e-13 b1=-4.033143240e-09 lb1=4.921294497e-14 pb1=2.646977960e-35 keta=-1.917560068e-02 lketa=8.548590692e-8 dwg=0.0 dwb=0.0 pclm=-3.426882576e-01 lpclm=3.389244816e-06 ppclm=1.332267630e-27 pdiblc1=0.39 pdiblc2=-1.025171335e-03 lpdiblc2=2.913057840e-8 pdiblcb=-0.025 drout=0.56 pscbe1=5.275926511e+08 lpscbe1=1.076521426e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.828274235e-01 lkt1=-1.223999366e-7 kt2=-1.864692104e-02 lkt2=-9.900092610e-8 at=1.698195537e+05 lat=-1.178433279e-1 ute=-8.085800536e-01 lute=-2.338011625e-6 ua1=2.387533168e-09 lua1=-7.149004768e-15 ub1=-1.684552764e-18 lub1=5.026803557e-24 uc1=-1.180400046e-11 luc1=2.510239413e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.165 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.063679854e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.411827189e-8 k1=5.224894914e-01 lk1=1.588745419e-7 k2=-2.118364742e-02 lk2=-7.475510716e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.115687121e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.716048642e-9 nfactor=2.711869382e+00 lnfactor=1.437815308e-6 eta0=0.08 etab=-0.07 u0=2.960672257e-02 lu0=7.891014271e-10 ua=-4.947617111e-10 lua=-4.594867802e-16 ub=1.352170129e-18 lub=3.594191158e-25 uc=-4.842565428e-12 luc=9.817486230e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.363604600e+04 lvsat=2.622624489e-1 a0=8.479396350e-01 la0=1.272744237e-6 ags=4.366510930e-01 lags=-3.284451492e-7 a1=0.0 a2=0.42385546 b0=4.869543535e-08 lb0=4.896208513e-14 b1=9.935730785e-09 lb1=-5.990382877e-15 keta=-1.264073531e-02 lketa=5.966089661e-08 pketa=-6.938893904e-30 dwg=0.0 dwb=0.0 pclm=-7.366646536e-01 lpclm=4.946192650e-06 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=-5.529034283e-04 lpdiblc2=2.726423184e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.057875285e-01 lkt1=-3.166433390e-8 kt2=-5.663636600e-02 lkt2=5.112883963e-8 at=140000.0 ute=-1.610417584e+00 lute=8.307548749e-7 ua1=-3.141532565e-10 lua1=3.527738482e-15 pua1=1.654361225e-36 ub1=5.536467272e-20 lub1=-1.849143105e-24 uc1=5.805098873e-11 luc1=-2.503466317e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.166 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.842615762e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.903080817e-8 k1=6.212681700e-01 lk1=-3.392968399e-8 k2=-6.424800454e-02 lk2=9.301393283e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.823954033e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.030090856e-8 nfactor=3.187048083e+00 lnfactor=5.103230289e-7 eta0=1.537410312e-01 leta0=-1.439337178e-7 etab=-1.363342072e-01 letab=1.294764787e-7 u0=3.391180834e-02 lu0=-7.613913680e-9 ua=-2.540776782e-10 lua=-9.292733711e-16 ub=1.172408749e-18 lub=7.102919370e-25 uc=4.822878123e-11 luc=-5.414090889e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.213473320e+05 lvsat=5.202283627e-2 a0=1.5 ags=3.313088529e-01 lags=-1.228296323e-7 a1=0.0 a2=0.42385546 b0=2.633747057e-07 lb0=-3.700663038e-13 b1=4.471577028e-09 lb1=4.674995022e-15 keta=1.805004733e-02 lketa=-2.438589030e-10 dwg=0.0 dwb=0.0 pclm=2.522733322e+00 lpclm=-1.415764330e-6 pdiblc1=2.001896837e-01 lpdiblc1=3.704871499e-7 pdiblc2=2.062764645e-02 lpdiblc2=-1.407768104e-8 pdiblcb=-0.025 drout=4.703102312e-01 ldrout=1.750637556e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.467909273e-01 lkt1=4.836942111e-8 kt2=-3.423300662e-02 lkt2=7.400148129e-9 at=1.495188100e+05 lat=-1.857958438e-2 ute=-1.628064281e+00 lute=8.651991289e-7 ua1=8.257868283e-10 lua1=1.302711089e-15 ub1=-4.438155885e-19 lub1=-8.748026374e-25 uc1=4.300065746e-11 luc1=4.341792472e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.167 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.871474887e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.628376289e-8 k1=5.947741785e-01 lk1=-8.710556888e-9 k2=-6.023609446e-02 lk2=5.482532296e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.191289451e-01 ldsub=3.890438058e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.073244113e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.165319250e-8 nfactor=3.993154312e+00 lnfactor=-2.569941745e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-1.387778781e-22 peta0=6.765421556e-29 etab=-0.0003125 u0=2.578130380e-02 lu0=1.253591093e-10 ua=-1.288073434e-09 lua=5.496754344e-17 ub=2.017358362e-18 lub=-9.399954564e-26 uc=7.700792919e-11 luc=-3.280841503e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.065995738e+05 lvsat=-2.912715290e-2 a0=1.5 ags=3.674223382e-01 lags=-1.572053728e-7 a1=0.0 a2=0.42385546 b0=-2.387298510e-07 lb0=1.078774838e-13 b1=1.786280847e-08 lb1=-8.071863754e-15 keta=3.545712353e-02 lketa=-1.681332400e-8 dwg=0.0 dwb=0.0 pclm=1.409768704e+00 lpclm=-3.563544566e-7 pdiblc1=6.704934226e-01 lpdiblc1=-7.718604331e-8 pdiblc2=9.917256884e-03 lpdiblc2=-3.882664709e-09 ppdiblc2=-3.469446952e-30 pdiblcb=-0.025 drout=3.417242576e-01 ldrout=2.974623007e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.851443400e-07 lalpha0=4.903561095e-13 walpha0=-1.058791184e-28 palpha0=2.646977960e-35 alpha1=0.85 beta0=1.228745412e+01 lbeta0=1.496876545e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.870790129e-01 lkt1=-8.469215655e-9 kt2=-5.289864105e-03 lkt2=-2.015027931e-8 at=2.474890600e+05 lat=-1.118356039e-1 ute=-2.741143519e-02 lute=-6.584319030e-7 ua1=3.835299287e-09 lua1=-1.561986640e-15 ub1=-2.642421110e-18 lub1=1.218008185e-24 uc1=-5.541599185e-12 luc1=5.054824427e-17 puc1=2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.168 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-4.948766302e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.600418038e-07 wvth0=4.437774325e-07 pvth0=-2.005345900e-13 k1=3.077427632e-01 lk1=1.209934861e-07 wk1=-6.000826502e-16 pk1=2.711657565e-22 k2=6.013024137e-02 lk2=-4.890872790e-08 wk2=-1.609685100e-08 pk2=7.273861128e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.920407444e+00 ldsub=-7.298710488e-07 wdsub=-7.327058495e-07 pdsub=3.310958520e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590366e-03 lcdscd=-1.221701118e-09 wcdscd=-5.447323148e-18 pcdscd=2.461541387e-24 cit=0.0 voff='-4.024725158e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.217186281e-07 wvoff=1.289225013e-07 pvoff=-5.825762879e-14 nfactor=-3.609281044e+00 lnfactor=3.178401917e-06 wnfactor=3.248580752e-06 pnfactor=-1.467971919e-12 eta0=8.778146603e-01 leta0=-1.752460369e-07 weta0=3.080560133e-09 peta0=-1.392046594e-15 etab=3.496458977e-02 letab=-1.594104660e-08 wetab=-2.591008961e-17 petab=1.170827432e-23 u0=-2.639517307e-02 lu0=2.370291766e-08 wu0=2.070304533e-08 pu0=-9.355312828e-15 ua=-1.029192944e-09 lua=-6.201563167e-17 wua=-5.539007474e-17 pua=2.502972236e-23 ub=2.677969457e-18 lub=-3.925171479e-25 wub=-4.864439007e-25 pub=2.198147563e-31 uc=-7.838167151e-11 luc=3.740919313e-17 wuc=4.886185059e-18 puc=-2.207974191e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.500141474e+05 lvsat=-3.557273836e-03 wvsat=-6.395088462e-03 pvsat=2.889818969e-9 a0=1.500000005e+00 la0=-2.116827602e-15 wa0=-1.833141638e-15 pa0=8.283613795e-22 ags=-9.741017959e-01 lags=4.490038944e-07 wags=-3.924924274e-16 pags=1.773598352e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.195796501e-01 lketa=-1.000147954e-07 wketa=-6.555742461e-08 pketa=2.962415459e-14 dwg=0.0 dwb=0.0 pclm=3.252942902e-01 lpclm=1.336989261e-07 wpclm=2.548271952e-07 ppclm=-1.151515678e-13 pdiblc1=6.149252007e-01 lpdiblc1=-5.207581962e-08 wpdiblc1=3.138298510e-16 ppdiblc1=-1.418136719e-22 pdiblc2=-4.393116251e-03 lpdiblc2=2.583921013e-09 wpdiblc2=-8.414493061e-18 ppdiblc2=3.802347760e-24 pdiblcb=3.822571344e-02 lpdiblcb=-2.857049861e-08 wpdiblcb=-2.491468143e-17 ppdiblcb=1.125849414e-23 drout=1.401075646e+00 ldrout=-1.812384642e-07 wdrout=-1.662172622e-15 pdrout=7.511045119e-22 pscbe1=8.069286532e+08 lpscbe1=-3.130926756e+00 wpscbe1=-1.642093658e-07 ppscbe1=7.420277596e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.383073786e-06 lalpha0=-3.538561654e-13 walpha0=-1.331385544e-13 palpha0=6.016278309e-20 alpha1=0.85 beta0=1.747630247e+01 lbeta0=-8.478654378e-07 wbeta0=-3.550361483e-07 pbeta0=1.604340897e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.475295498e-01 lkt1=-7.152896660e-08 wkt1=-8.875903695e-08 pkt1=4.010852237e-14 kt2=-6.684223721e-02 lkt2=7.664068600e-09 wkt2=-9.960088310e-18 pkt2=4.500788631e-24 at=1.348084708e+05 lat=-6.091738660e-02 wat=-6.656927767e-02 pat=3.008139176e-8 ute=-1.196779523e+00 lute=-1.300166823e-07 wute=-1.775180737e-07 pute=8.021704467e-14 ua1=7.037062504e-10 lua1=-1.468792468e-16 wua1=-1.879303894e-24 pua1=8.492215638e-31 ub1=-4.757344990e-19 lub1=2.389236724e-25 wub1=-2.669641274e-33 pub1=1.206360111e-39 uc1=7.331997412e-11 luc1=1.491219767e-17 wuc1=3.865456361e-26 puc1=-1.746726280e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.169 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.429716875e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.341400576e-07 wvth0=-1.584919402e-06 pvth0=2.090207556e-13 k1=9.070734845e-01 lk1=7.222720200e-16 wk1=2.143149658e-15 pk1=-2.826407997e-22 k2=-2.781048764e-01 lk2=1.937451590e-08 wk2=5.748875358e-08 pk2=-7.581674311e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-6.063362996e+00 ldsub=8.819005114e-07 wdsub=2.616806605e-06 pdsub=-3.451070719e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999950e-03 lcdscd=6.556510543e-18 wcdscd=1.945470868e-17 pcdscd=-2.565706328e-24 cit=0.0 voff='9.690905439e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.551738940e-07 wvoff=-4.604375045e-07 pvoff=6.072295853e-14 nfactor=3.150280748e+01 lnfactor=-3.910061627e-06 wnfactor=-1.160207411e-05 pnfactor=1.530093136e-12 eta0=2.811495795e-02 leta0=-3.707828399e-09 weta0=-1.100200048e-08 peta0=1.450954825e-15 etab=-4.399800024e-02 letab=3.118591496e-17 wetab=9.253597888e-17 petab=-1.220373802e-23 u0=2.144474425e-01 lu0=-2.491863041e-08 wu0=-7.393944761e-08 pu0=9.751208291e-15 ua=-1.666619528e-09 lua=6.666868467e-17 wua=1.978216955e-16 pua=-2.608892302e-23 ub=-2.166525487e-18 lub=5.854943359e-25 wub=1.737299645e-24 pub=-2.291168145e-31 uc=1.360531218e-10 luc=-5.881117375e-18 wuc=-1.745066093e-17 puc=2.301410613e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.426576204e+04 lvsat=7.697265947e-03 wvsat=2.283960165e-02 pvsat=-3.012109505e-9 a0=1.499999983e+00 la0=2.206405725e-15 wa0=6.546930109e-15 pa0=-8.634155613e-22 ags=1.249999996e+00 lags=4.724123315e-16 wags=1.401758709e-15 pags=-1.848654563e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.666905832e-01 lketa=7.890632554e-08 wketa=2.341336593e-07 pketa=-3.087778112e-14 dwg=0.0 dwb=0.0 pclm=2.506848851e+00 lpclm=-3.067154901e-07 wpclm=-9.100971256e-07 ppclm=1.200245190e-13 pdiblc1=3.569721529e-01 lpdiblc1=-3.777322899e-16 wpdiblc1=-1.120820770e-15 ppdiblc1=1.478149825e-22 pdiblc2=8.406112023e-03 lpdiblc2=1.012785689e-17 wpdiblc2=3.005176663e-17 ppdiblc2=-3.963253337e-24 pdiblcb=-1.032957702e-01 lpdiblcb=2.998790105e-17 wpdiblcb=8.898104475e-17 ppdiblcb=-1.173491859e-23 drout=5.033266448e-01 ldrout=2.000627219e-15 wdrout=5.936332315e-15 pdrout=-7.828893089e-22 pscbe1=7.914198785e+08 lpscbe1=1.976451874e-07 wpscbe1=5.864601135e-07 ppscbe1=-7.734298706e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.163498658e-06 lalpha0=1.602484261e-13 walpha0=4.754948371e-13 palpha0=-6.270873461e-20 alpha1=0.85 beta0=1.115973688e+01 lbeta0=4.273291403e-07 wbeta0=1.267986244e-06 pbeta0=-1.672232938e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.031026518e+00 lkt1=1.068322849e-07 wkt1=3.169965605e-07 pkt1=-4.180582340e-14 kt2=-2.887893909e-02 lkt2=1.198821598e-17 wkt2=3.557182326e-17 pkt2=-4.691247391e-24 at=-5.638288464e+05 lat=8.012421364e-02 wat=2.377474203e-01 pat=-3.135436753e-8 ute=-2.899174755e+00 lute=2.136645696e-07 wute=6.339931204e-07 pute=-8.361164671e-14 ua1=-2.384735315e-11 lua1=2.261970104e-24 wua1=6.711798291e-24 pua1=-8.851586710e-31 ub1=7.077531456e-19 lub1=3.213237697e-33 wub1=9.534433286e-33 pub1=-1.257410387e-39 uc1=1.471862504e-10 luc1=-4.652549734e-26 wuc1=-1.380518947e-25 puc1=1.820645208e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.170 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-2.522595364e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.827378328e-07 wvth0=1.366349450e-06 pvth0=-1.801955318e-13 k1=0.90707349 k2=-1.214234996e+00 lk2=1.428322922e-07 wk2=4.202331718e-07 pk2=-5.542077093e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.091390987e+00 ldsub=-3.254375986e-07 wdsub=-1.039679862e-06 pdsub=1.371140199e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-5.755837948e+00 lnfactor=1.003645791e-06 wnfactor=2.035947004e-06 pnfactor=-2.685027268e-13 eta0=3.773678949e-04 leta0=-4.976765037e-11 weta0=-1.589933803e-10 peta0=2.096820599e-17 etab=-0.043998 u0=1.180195927e-01 lu0=-1.220162915e-08 wu0=-3.513079141e-08 pu0=4.633083902e-15 ua=-1.561180192e-09 lua=5.276323956e-17 wua=2.136372329e-16 pua=-2.817469192e-23 ub=3.405756539e-18 lub=-1.493837899e-25 wub=-2.026061243e-25 pub=2.671989827e-32 uc=-1.174583905e-10 luc=2.755223438e-17 wuc=1.212251842e-16 puc=-1.598729852e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.803855899e+05 lvsat=-5.641270307e-02 wvsat=-1.776827075e-01 pvsat=2.343297315e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-9.287045780e-01 lketa=1.134609932e-07 wketa=3.968494623e-07 pketa=-5.233690393e-14 dwg=0.0 dwb=0.0 pclm=2.580727704e-02 lpclm=2.048675365e-08 wpclm=1.189334913e-07 ppclm=-1.568506776e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.249543128e-07 lalpha0=-9.674040130e-15 walpha0=3.020736542e-21 palpha0=-3.983777534e-28 alpha1=0.85 beta0=1.626781828e+01 lbeta0=-2.463297431e-07 wbeta0=2.089785767e-14 pbeta0=-2.756024742e-21 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.530400709e-01 lkt1=-8.957445766e-09 wkt1=-1.040710629e-15 pkt1=1.372498781e-22 kt2=-0.028878939 at=9.760154460e+03 lat=4.478722616e-03 wat=-3.342397977e-10 pat=4.407987581e-17 ute=-9.447486384e-01 lute=-4.408710108e-08 wute=-2.266950667e-07 pute=2.989677209e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.171 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.4922131+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.039695546 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.8826 eta0=0.08 etab=-0.07 u0=0.0266513 ua=-1.0573461e-9 ub=1.802952e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=6.3469e-8 b1=2.5194e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.172 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.814679883e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.143851906e-7 k1=5.567098995e-01 lk1=2.254127697e-7 k2=-3.239100444e-02 lk2=-1.457393440e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017808550e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.296270710e-7 nfactor=2.951582568e+00 lnfactor=-1.376331981e-6 eta0=0.08 etab=-0.07 u0=2.560927226e-02 lu0=2.079041345e-8 ua=-1.145242396e-09 lua=1.753696429e-15 ub=1.844100334e-18 lub=-8.209866543e-25 uc=6.327183549e-11 luc=-2.939876843e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.478299869e+00 la0=-2.308430009e-6 ags=3.215147230e-01 lags=4.661812263e-7 a1=0.0 a2=0.42385546 b0=5.268624936e-08 lb0=2.151361575e-13 b1=2.760408260e-09 lb1=-4.808568123e-15 keta=-1.976419529e-03 lketa=-5.127993490e-8 dwg=0.0 dwb=0.0 pclm=-2.729504833e-02 lpclm=8.812755480e-07 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=-1.515165620e-04 lpdiblc2=2.218337962e-08 ppdiblc2=-6.938893904e-30 pdiblcb=-0.025 drout=0.56 pscbe1=-6.522518163e+07 lpscbe1=5.790538287e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.785341441e-01 lkt1=-1.565395837e-7 kt2=-2.847160196e-02 lkt2=-2.087623258e-08 wkt2=-2.775557562e-23 at=1.882531350e+05 lat=-2.644249724e-1 ute=-1.123882006e+00 lute=1.692319823e-7 ua1=8.774736444e-10 lua1=4.858808868e-15 ub1=-2.494531757e-19 lub1=-6.384937596e-24 uc1=4.313166665e-11 luc1=-1.858179462e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.173 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.164933975e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-6.413269591e-8 k1=6.071532016e-01 lk1=-1.757063659e-7 k2=-6.120959896e-02 lk2=8.342269022e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.259465233e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.253544744e-8 nfactor=2.484875242e+00 lnfactor=2.334869137e-6 eta0=0.08 etab=-0.07 u0=2.666023828e-02 lu0=1.243325671e-8 ua=-1.234602158e-09 lua=2.464274623e-15 ub=2.035011298e-18 lub=-2.339087928e-24 uc=3.252620055e-11 luc=-4.950205394e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.205783465e+00 la0=-1.414119935e-7 ags=4.064200086e-01 lags=-2.089755015e-7 a1=0.0 a2=0.42385546 b0=9.817257298e-08 lb0=-1.465656750e-13 b1=-4.033143240e-09 lb1=4.921294497e-14 keta=-1.917560068e-02 lketa=8.548590692e-8 dwg=0.0 dwb=0.0 pclm=-3.426882576e-01 lpclm=3.389244816e-06 wpclm=-1.110223025e-22 pdiblc1=0.39 pdiblc2=-1.025171335e-03 lpdiblc2=2.913057840e-08 ppdiblc2=-1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=5.275926511e+08 lpscbe1=1.076521426e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.828274235e-01 lkt1=-1.223999366e-7 kt2=-1.864692104e-02 lkt2=-9.900092610e-8 at=1.698195537e+05 lat=-1.178433279e-1 ute=-8.085800536e-01 lute=-2.338011625e-6 ua1=2.387533168e-09 lua1=-7.149004768e-15 pua1=6.617444900e-36 ub1=-1.684552764e-18 lub1=5.026803557e-24 uc1=-1.180400046e-11 luc1=2.510239413e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.174 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='5.063679854e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.411827189e-8 k1=5.224894914e-01 lk1=1.588745419e-7 k2=-2.118364742e-02 lk2=-7.475510716e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.115687121e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.716048642e-9 nfactor=2.711869382e+00 lnfactor=1.437815308e-6 eta0=0.08 etab=-0.07 u0=2.960672257e-02 lu0=7.891014271e-10 ua=-4.947617111e-10 lua=-4.594867802e-16 ub=1.352170129e-18 lub=3.594191158e-25 uc=-4.842565428e-12 luc=9.817486230e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.363604600e+04 lvsat=2.622624489e-1 a0=8.479396350e-01 la0=1.272744237e-6 ags=4.366510930e-01 lags=-3.284451492e-7 a1=0.0 a2=0.42385546 b0=4.869543535e-08 lb0=4.896208513e-14 b1=9.935730785e-09 lb1=-5.990382877e-15 keta=-1.264073531e-02 lketa=5.966089661e-08 wketa=-3.469446952e-24 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=-7.366646536e-01 lpclm=4.946192650e-06 ppclm=1.776356839e-27 pdiblc1=0.39 pdiblc2=-5.529034283e-04 lpdiblc2=2.726423184e-08 ppdiblc2=-1.387778781e-29 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.057875285e-01 lkt1=-3.166433390e-8 kt2=-5.663636600e-02 lkt2=5.112883963e-8 at=140000.0 ute=-1.610417584e+00 lute=8.307548749e-7 ua1=-3.141532565e-10 lua1=3.527738482e-15 pua1=1.654361225e-36 ub1=5.536467272e-20 lub1=-1.849143105e-24 uc1=5.805098873e-11 luc1=-2.503466317e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.175 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.842615762e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.903080817e-8 k1=6.212681700e-01 lk1=-3.392968399e-8 k2=-6.424800454e-02 lk2=9.301393283e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.455643000e-01 ldsub=-5.573875314e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.823954033e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.030090856e-8 nfactor=3.187048083e+00 lnfactor=5.103230289e-7 eta0=1.537410312e-01 leta0=-1.439337178e-7 etab=-1.363342072e-01 letab=1.294764787e-7 u0=3.391180834e-02 lu0=-7.613913680e-9 ua=-2.540776782e-10 lua=-9.292733711e-16 ub=1.172408749e-18 lub=7.102919370e-25 uc=4.822878123e-11 luc=-5.414090889e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.213473320e+05 lvsat=5.202283627e-2 a0=1.5 ags=3.313088529e-01 lags=-1.228296323e-7 a1=0.0 a2=0.42385546 b0=2.633747057e-07 lb0=-3.700663038e-13 wb0=1.058791184e-28 pb0=1.058791184e-34 b1=4.471577028e-09 lb1=4.674995022e-15 keta=1.805004733e-02 lketa=-2.438589030e-10 dwg=0.0 dwb=0.0 pclm=2.522733322e+00 lpclm=-1.415764330e-6 pdiblc1=2.001896837e-01 lpdiblc1=3.704871499e-7 pdiblc2=2.062764645e-02 lpdiblc2=-1.407768104e-8 pdiblcb=-0.025 drout=4.703102312e-01 ldrout=1.750637556e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.467909273e-01 lkt1=4.836942111e-8 kt2=-3.423300662e-02 lkt2=7.400148129e-9 at=1.495188100e+05 lat=-1.857958438e-2 ute=-1.628064281e+00 lute=8.651991289e-7 ua1=8.257868283e-10 lua1=1.302711089e-15 ub1=-4.438155885e-19 lub1=-8.748026374e-25 uc1=4.300065746e-11 luc1=4.341792472e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.176 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='4.871474887e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.628376289e-8 k1=5.947741785e-01 lk1=-8.710556888e-9 k2=-6.023609446e-02 lk2=5.482532296e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.191289451e-01 ldsub=3.890438058e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.073244113e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.165319250e-8 nfactor=3.993154312e+00 lnfactor=-2.569941745e-7 eta0=-4.380244824e-01 leta0=4.193566311e-07 weta0=-1.734723476e-23 peta0=-1.006139616e-28 etab=-0.0003125 u0=2.578130380e-02 lu0=1.253591093e-10 ua=-1.288073434e-09 lua=5.496754344e-17 ub=2.017358362e-18 lub=-9.399954564e-26 uc=7.700792919e-11 luc=-3.280841503e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.065995738e+05 lvsat=-2.912715290e-2 a0=1.5 ags=3.674223382e-01 lags=-1.572053728e-7 a1=0.0 a2=0.42385546 b0=-2.387298510e-07 lb0=1.078774838e-13 b1=1.786280847e-08 lb1=-8.071863754e-15 keta=3.545712353e-02 lketa=-1.681332400e-8 dwg=0.0 dwb=0.0 pclm=1.409768704e+00 lpclm=-3.563544566e-7 pdiblc1=6.704934226e-01 lpdiblc1=-7.718604331e-8 pdiblc2=9.917256884e-03 lpdiblc2=-3.882664709e-09 wpdiblc2=6.938893904e-24 pdiblcb=-0.025 drout=3.417242576e-01 ldrout=2.974623007e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-4.851443400e-07 lalpha0=4.903561095e-13 walpha0=1.588186776e-28 palpha0=5.293955920e-35 alpha1=0.85 beta0=1.228745412e+01 lbeta0=1.496876545e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-2.870790129e-01 lkt1=-8.469215655e-9 kt2=-5.289864105e-03 lkt2=-2.015027931e-8 at=2.474890600e+05 lat=-1.118356039e-1 ute=-2.741143519e-02 lute=-6.584319030e-7 ua1=3.835299287e-09 lua1=-1.561986640e-15 ub1=-2.642421110e-18 lub1=1.218008185e-24 uc1=-5.541599185e-12 luc1=5.054824427e-17 puc1=2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.177 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='6.391700947e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.241236434e-8 k1=3.077427617e-01 lk1=1.209934868e-7 k2=1.899569999e-02 lk2=-3.032081021e-08 pk2=1.387778781e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.802140521e-02 ldsub=1.162246268e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.103590352e-03 lcdscd=-1.221701112e-09 wcdscd=-6.938893904e-24 cit=0.0 voff='-7.301876348e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.715526294e-8 nfactor=4.692273051e+00 lnfactor=-5.729126495e-7 eta0=8.856867600e-01 leta0=-1.788033288e-7 etab=3.496458970e-02 letab=-1.594104657e-08 wetab=1.734723476e-24 petab=1.626303259e-30 u0=2.651022282e-02 lu0=-2.040255453e-10 ua=-1.170738972e-09 lua=1.946328970e-18 ub=1.434891121e-18 lub=1.692063338e-25 uc=-6.589531741e-11 luc=3.176684695e-17 wuc=6.462348536e-33 puc=9.693522803e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.336718808e+05 lvsat=3.827485950e-3 a0=1.5 ags=-9.741017969e-01 lags=4.490038949e-07 wags=-3.053113318e-22 pags=-8.326672685e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.205156677e-02 lketa=-2.431203761e-08 wketa=-3.469446952e-24 pketa=-4.770489559e-30 dwg=0.0 dwb=0.0 pclm=9.764899684e-01 lpclm=-1.605640282e-7 pdiblc1=6.149252015e-01 lpdiblc1=-5.207581998e-8 pdiblc2=-4.393116272e-03 lpdiblc2=2.583921023e-9 pdiblcb=3.822571337e-02 lpdiblcb=-2.857049858e-08 ppdiblcb=1.387778781e-29 drout=1.401075642e+00 ldrout=-1.812384623e-7 pscbe1=8.069286528e+08 lpscbe1=-3.130926566e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.042846162e-06 lalpha0=-2.001137663e-13 alpha1=0.85 beta0=1.656902880e+01 lbeta0=-4.378857032e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-3.743479677e-01 lkt1=3.096596692e-8 kt2=-6.684223724e-02 lkt2=7.664068612e-9 at=-3.530534254e+04 lat=1.595381349e-2 ute=-1.650416358e+00 lute=7.497318452e-8 ua1=7.037062456e-10 lua1=-1.468792446e-16 ub1=-4.757345058e-19 lub1=2.389236755e-25 wub1=9.629649722e-41 pub1=-7.222237291e-47 uc1=7.331997422e-11 luc1=1.491219762e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.178 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='0.37955+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.90707349 k2=-0.1311958 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.62373 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=1.8544 eta0=0.0 etab=-0.043998 u0=0.0254996 ua=-1.161098e-9 ub=2.27304e-18 uc=9.1459e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=152631.0 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.068376 dwg=0.0 dwb=0.0 pclm=0.18115 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.16e-8 alpha1=0.85 beta0=14.4 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=43720.487 ute=-1.2790432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.179 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='3.996598e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.9635*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=-6.60999999999998e-10 lint=2.40595e-8 vth0='-3.719569900e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.910949335e-08 wvth0=5.247573396e-07 pvth0=-6.920552270e-14 k1=0.90707349 k2=-4.158704441e-01 lk2=3.754317674e-08 wk2=1.078155588e-07 pk2=-1.421882371e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.145270833e+00 ldsub=-3.325433265e-07 wdsub=-1.060764231e-06 pdsub=1.398946476e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-5.755837763e+00 lnfactor=1.003645766e-06 wnfactor=2.035946931e-06 pnfactor=-2.685027173e-13 eta0=6.038887884e-04 leta0=-7.964144934e-11 weta0=-2.476359805e-10 peta0=3.265848075e-17 etab=-0.043998 u0=2.605260337e-02 lu0=-7.293063698e-11 wu0=8.579147789e-10 pu0=-1.131426590e-16 ua=-1.561180684e-09 lua=5.276330447e-17 wua=2.136374256e-16 pua=-2.817471732e-23 ub=3.405791239e-18 lub=-1.493883661e-25 wub=-2.026197031e-25 pub=2.672168906e-32 uc=-1.237407073e-10 luc=2.838075260e-17 wuc=1.236835930e-16 puc=-1.631151593e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.566624309e+05 lvsat=-1.371976914e-02 wvsat=-5.100271349e-02 pvsat=6.726288858e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-9.287047565e-01 lketa=1.134610167e-07 wketa=3.968495321e-07 pketa=-5.233691314e-14 dwg=0.0 dwb=0.0 pclm=2.580720676e-02 lpclm=2.048676292e-08 wpclm=1.189335188e-07 ppclm=-1.568507139e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.249543200e-07 lalpha0=-9.674041071e-15 walpha0=2.285430417e-22 palpha0=-3.014048952e-29 alpha1=0.85 beta0=1.626781834e+01 lbeta0=-2.463297501e-07 wbeta0=4.001776688e-17 pbeta0=-5.275779813e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=1.85814e-8 dwc=-2.252e-8 xpart=0.0 cgso=2.4133302e-10 cgdo=2.4133302e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001131080901 mjs=0.44 pbsws=0.2 cjsws=3.101378147e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.011274009e-10 mjswgs=0.8 tnom=30.0 kt1=-1.530400733e-01 lkt1=-8.957445444e-09 wkt1=-8.505551818e-17 pkt1=1.121713833e-23 kt2=-0.028878939 at=9.760153675e+03 lat=4.478722719e-03 wat=-2.698588651e-11 pat=3.558932804e-18 ute=-9.330005132e-01 lute=-4.563645557e-08 wute=-2.312923665e-07 pute=3.050306858e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.ends sky130_fd_pr__nfet_01v8