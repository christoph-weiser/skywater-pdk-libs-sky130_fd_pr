* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8_lvt__toxe_mult=0.948
.param sky130_fd_pr__nfet_01v8_lvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__overlap_mult=0.86067
.param sky130_fd_pr__nfet_01v8_lvt__ajunction_mult=0.82447
.param sky130_fd_pr__nfet_01v8_lvt__pjunction_mult=0.75
.param sky130_fd_pr__nfet_01v8_lvt__lint_diff=1.7325e-8
.param sky130_fd_pr__nfet_01v8_lvt__wint_diff=-3.2175e-8
.param sky130_fd_pr__nfet_01v8_lvt__dlc_diff=1.1336e-8
.param sky130_fd_pr__nfet_01v8_lvt__dwc_diff=-3.2175e-8
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_0=-0.10724
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_0=-0.093222
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_0=0.0081846
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_0=0.0013057
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0=0.0023529
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_0=-0.1697
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_0=2.7218e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_0=3.8431e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0=0.30318
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0=-0.0046766
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_1=-0.072473
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_1=-0.096311
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_1=0.0080507
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1=0.00147426
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_1=-0.14919
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_1=0.00011578
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_1=2.8356e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_1=2.6855e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1=0.27456
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1=-0.0063307
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2=-0.00037846
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_2=0.0046126
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_2=-0.11674
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_2=0.010192
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2=0.001
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_2=-0.019102
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_2=-6.7162e-5
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_2=-4.0716e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_2=2.4704e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2=0.30957
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3=-0.12083
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3=0.071167
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3=-0.06459
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_3=-0.024322
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_3=0.0504
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3=0.0045
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_3=-0.0025347
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_3=2.99e-11
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3=-37719.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_3=1.9717e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4=-0.044924
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4=0.18285
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4=-0.067816
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_4=-0.077947
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_4=0.030667
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4=0.0035327
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_4=-0.0027063
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_4=1.4975e-11
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4=-27268.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_4=9.1673e-20
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_5=4.9257e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5=0.38483
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5=-0.0077756
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_5=-0.11254
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_5=0.012134
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5=0.0010833
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_5=0.00182
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_5=1.0925e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5=-18670.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_6=2.7039e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6=0.33805
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6=-0.0062083
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_6=-0.10389
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_6=-0.0011301
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6=0.0030639
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_6=-0.00026232
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_6=-1.4498e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6=-16312.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_7=2.237e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7=0.24768
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7=0.0049372
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_7=-0.044883
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_7=-0.083842
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_7=0.0033279
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7=0.0016389
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_7=-0.052674
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_7=0.00077332
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_7=-3.0348e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8=0.00199938
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_8=-0.051192
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_8=8.7555e-5
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_8=9.4746e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_8=1.7506e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8=0.2391
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8=-0.0028836
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_8=-0.03459
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_8=-0.086594
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_8=0.00064808
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9=0.0021675
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_9=-0.017152
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_9=-0.00027835
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_9=-1.8365e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_9=1.1976e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9=0.23485
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9=0.0031712
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_9=0.0040339
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_9=-0.09247
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_9=0.0056151
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_10=2.6243e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_10=-1.4198e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10=0.0031233
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_10=-0.0046344
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10=-30297.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10=-0.067091
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10=-0.73159
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10=-0.083472
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_10=0.0045616
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_10=0.054313
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_11=0.033481
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_11=1.9818e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_11=9.3123e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11=0.0036808
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_11=-0.0019243
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11=-19197.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11=-0.03687
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11=0.29166
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11=-0.041779
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_11=-0.094472
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_12=0.02058
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_12=1.2994e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_12=3.7224e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12=0.00083124
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_12=0.00095499
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12=-9309.5
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12=-0.0026687
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12=0.41021
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_12=-0.11654
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_13=0.012552
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_13=1.7628e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_13=2.2271e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13=0.0015175
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_13=-0.00041587
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13=-7419.7
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13=0.0038312
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13=0.29916
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_13=-0.095191
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14=0.22224
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_14=-0.073593
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_14=0.002812
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_14=9.5412e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_14=1.9897e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_14=-0.05226
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14=0.00197129
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_14=-0.071021
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_14=0.00038113
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14=-0.0045428
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15=0.0053271
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15=0.22251
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_15=-0.085479
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_15=-0.0061278
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_15=-5.7198e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_15=2.1734e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_15=0.0029657
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15=0.002009
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_15=0.0048954
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_15=0.0004302
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16=0.0018021
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_16=-0.03219
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_16=-2.8938e-5
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16=-0.0095281
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16=0.20081
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_16=-0.078124
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_16=0.0081435
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_16=1.1846e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_16=1.4143e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_16=0.0045892
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17=0.0035038
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_17=-0.0026687
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17=-26507.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17=-0.074112
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17=-0.052134
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_17=-0.0013863
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_17=0.057166
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_17=3.0202e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_17=6.2924e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18=0.0013916
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_18=-0.0024675
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18=-22692.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18=-0.022761
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18=0.15638
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_18=-0.051155
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_18=0.03356
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_18=1.2859e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_18=5.063e-20
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_19=3.0062e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19=0.0017707
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_19=-0.00019199
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19=-15177.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19=-0.012464
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19=0.34467
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_19=-0.094448
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_19=0.013596
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_19=3.5652e-12
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_20=-3.9165e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_20=2.3083e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20=0.0016075
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_20=0.00010669
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20=-3727.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20=-0.0012631
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20=0.27695
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_20=-0.088637
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_20=0.0015349
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_21=-2.5325e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_21=2.2719e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_21=0.036717
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21=0.0014
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_21=0.043576
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_21=0.00081759
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21=0.0059539
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21=0.2405
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_21=-0.091068
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_21=-0.0052929
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_22=0.007281
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_22=4.94e-15
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_22=1.709e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_22=-0.0071609
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22=0.002
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_22=-0.01746
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_22=0.00018433
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22=-0.00251
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22=0.20821
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_22=-0.077032
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_23=0.0064536
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_23=-1.5075e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_23=1.907e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_23=-0.0024648
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23=-0.0004
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_23=0.022769
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_23=0.0005228
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23=-0.0027939
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23=0.25136
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23=-0.1
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_23=-0.1032
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_24=0.05951
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_24=4.032e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_24=-2.4003e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24=0.0010928
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_24=-0.005
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24=-24843.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24=-0.030521
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24=-1.5
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_24=-0.039992
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25=0.2288
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_25=-0.065769
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_25=0.032673
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_25=1.2484e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_25=-2.7509e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25=0.002603
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_25=-0.0028902
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25=-17841.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25=-0.020508
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26=-0.0088834
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26=0.32002
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_26=-0.089896
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_26=0.015591
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_26=2.3711e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_26=3.4661e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26=0.0010535
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_26=0.00065281
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26=-14474.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27=0.0014074
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_27=1.2597e-6
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27=-3404.1
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27=0.00246
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27=0.25902
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_27=-0.082883
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_27=0.0037121
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_27=-1.3023e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_27=1.9461e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28=0.0012
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_28=0.0013082
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28=-0.024114
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28=0.25608
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_28=-0.080102
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_28=1.8999e-7
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_28=1.1506e-8
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_28=0.0065995
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_28=2.1038e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_28=5.2387e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29=0.0041602
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_29=-0.0024166
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29=-36771.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29=-0.10687
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29=-0.060066
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29=-0.024775
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_29=-0.063748
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_29=0.04922
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_29=4.2051e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_29=2.7257e-19
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_30=7.8237e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30=0.0015098
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_30=-0.002199
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30=-35936.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30=-0.11916
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30=0.074462
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_30=-0.061736
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_30=0.021285
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_30=3.7522e-11
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_31=9.4623e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_31=-3.1689e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31=0.0044313
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_31=-0.0028421
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31=-43027.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31=-0.11958
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31=-0.068776
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31=-0.071833
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_31=-0.047169
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_31=0.032738
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_32=2.3172e-10
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_32=-4.2095e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32=0.0038442
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_32=-0.00067444
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32=-31335.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32=-0.13172
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32=-0.2
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32=-0.086428
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_32=-0.011311
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_32=0.033141
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_33=0.032169
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_33=8.1829e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_33=-2.9805e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33=0.0044325
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_33=-0.0018325
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33=-23311.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33=-0.11599
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33=-0.048661
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33=-0.07335
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_33=-0.044428
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_34=0.073427
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_34=1.061e-10
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_34=-3.9012e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34=0.0032691
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_34=-0.005
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34=-37559.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34=-0.06268
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34=-1.5
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34=-0.071509
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_34=-0.013658
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_35=0.07411
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_35=1.2347e-10
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_35=-3.0793e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35=0.0031992
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_35=-0.0046648
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35=-31504.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35=-0.064375
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35=-0.66492
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35=-0.084604
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_35=0.0035949
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36=0.052626
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_36=-0.020055
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_36=0.077414
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_36=6.5275e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_36=-8.7238e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36=0.0018875
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_36=-0.0036229
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36=-25852.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36=-0.068536
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37=-0.011492
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37=0.36824
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_37=-0.097534
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_37=0.027159
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_37=2.7122e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_37=-3.3913e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37=0.0018455
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_37=-0.0032585
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37=-13782.0
.include "sky130_fd_pr__nfet_01v8_lvt.pm3.spice"