* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__ind_05_220 a b ct sub
r31 net27 b r='1e-2'
r26 a net23 r='1e-2'
c2 net27 net31 c='223.7e-15'
c24 net35 net27 c='205e-15'
c25 net23 net37 c='223.7e-15'
r5 sub net31 r='5.358e3'
r4 net41 net27 r='2.059'
r13 net23 net35 r='9.064'
r10 sub net37 r='5.358e3'
r9 net23 net39 r='2.059'
l1 net39 ct l=4.96e-9
l3 ct net41 l=4.96e-9
.ends sky130_fd_pr__ind_05_220