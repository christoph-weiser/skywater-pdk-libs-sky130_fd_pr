* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre=0.0
.param sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre=0.0
.param sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre=0.0
.subckt sky130_fd_pr__rf_nfet_01v8_bm02 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_01v8_bm02 d g s b sky130_fd_pr__rf_nfet_01v8_bm02__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.0 nmos lmin=1.45e-07 lmax=1.55e-07 wmin=1.645e-06 wmax=1.655e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.90 rnoib=0.36 tnoia=2.7e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.633+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_0+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_0' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_0' ua='-1.96e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_0' ub='2.15e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_0' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_0' prwb=0.008 prwg=0.0 wr=1.0 u0='0.036+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_0' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_0' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_0' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_0' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_0' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.206+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_0+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='2.808+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_0' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.3121 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.2481 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.290+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_0' kt2=-0.02437 at=5.978e+4 ute=-1.681 ua1=6.012e-10 ub1=-4.98e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='900*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='7.7e-07+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.659e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.84e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='1e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.58e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='4.21e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.1 nmos lmin=1.75e-07 lmax=1.85e-07 wmin=1.645e-06 wmax=1.655e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-5.408e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.90 rnoib=0.36 tnoia=2.7e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.6345+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_1+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_1' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_1' ua='-1.985e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_1' ub='2.161e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_1' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_1' prwb=0.008 prwg=0.0 wr=1.0 u0='0.037+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_1' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_1' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_1' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_1' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_1' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1854+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_1+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.629+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_1' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.3121 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.2293 pdiblc2=0.016 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.02336 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2779+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_1' kt2=-0.02437 at=6.122e+4 ute=-1.5633 ua1=6.012e-10 ub1=-6.52e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='900*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.12e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.0 tpbsw=0.0 tpbswg=0.0 tcj=0.000992 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.629e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='4e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='1e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.18e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.41e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.2 nmos lmin=2.45e-07 lmax=2.55e-07 wmin=1.645e-06 wmax=1.655e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-5.408e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.90 rnoib=0.36 tnoia=2.7e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.625+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_2+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_2' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.564e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_2' ua='-1.985e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_2' ub='2.202e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_2' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_2' prwb=0.008 prwg=0.0 wr=1.0 u0='0.031+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_2' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_2' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_2' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_2' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_2' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1854+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_2+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.629+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_2' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.3121 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.04127 pdiblc2=0.01376 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.02336 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2779+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_2' kt2=-0.02437 at=5.449e+4 ute=-1.5633 ua1=6.012e-10 ub1=-6.52e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='900*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.35e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.629e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='4.1e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='1e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='8e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='1.7e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.41e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.ends sky130_fd_pr__rf_nfet_01v8_bm02
.subckt sky130_fd_pr__rf_nfet_01v8_bm02w3p00 d g s b
.param l=1
.param w=3.01
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_01v8_bm02w3p00 d g s b sky130_fd_pr__rf_nfet_01v8_bm02__model l='l' w=3.01 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.3 nmos lmin=1.45e-07 lmax=1.55e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.59+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_3+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_3' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_3' ua='-2.032e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_3' ub='2.05e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_3' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_3' prwb=0.008 prwg=0.0 wr=1.0 u0='0.03599+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_3' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_3' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_3' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_3' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_3' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1943+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_3+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='3.052+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_3' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.5779 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.2481 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.290+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_3' kt2=-0.02437 at=6.698e+4 ute=-1.5297 ua1=6.012e-10 ub1=-3.37e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='440*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='8.6e-07+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.0 tpbsw=0.0 tpbswg=0.0 tcj=0.000992 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.489e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.7e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.58e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.01e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.4 nmos lmin=1.75e-07 lmax=1.85e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.618+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_4+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_4' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.57e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_4' ua='-2.032e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_4' ub='2.124e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_4' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_4' prwb=0.008 prwg=0.0 wr=1.0 u0='0.03199+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_4' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_4' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_4' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_4' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_4' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1943+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_4+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.8+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_4' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.5779 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.1768 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03138 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.290+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_4' kt2=-0.02437 at=6.698e+4 ute=-1.5297 ua1=6.012e-10 ub1=-3.37e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='440*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.489e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.5e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.68e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.01e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.15 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.5 nmos lmin=2.45e-07 lmax=2.55e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.605+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_5+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_5' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.475e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_5' ua='-2.046e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_5' ub='2.28e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_5' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_5' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0275+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_5' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_5' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_5' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_5' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_5' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1943+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_5+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.8+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_5' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.5779 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.1768 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03138 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.290+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_5' kt2=-0.02437 at=6.698e+4 ute=-1.5297 ua1=6.012e-10 ub1=-3.37e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='440*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.35e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.889e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.6e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.68e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.71e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.15 pbswgs=0.9064
.ends sky130_fd_pr__rf_nfet_01v8_bm02w3p00
.subckt sky130_fd_pr__rf_nfet_01v8_bm02w5p00 d g s b
.param l=1
.param w=5.05
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_01v8_bm02w5p00 d g s b sky130_fd_pr__rf_nfet_01v8_bm02__model l='l' w=5.05 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.6 nmos lmin=1.45e-07 lmax=1.55e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.773e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.59+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_6+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_6' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_6' ua='-2.032e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_6' ub='2.12e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_6' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_6' prwb=0.008 prwg=0.0 wr=1.0 u0='0.03599+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_6' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_6' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_6' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_6' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_6' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1943+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_6+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='3.052+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_6' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.4128 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.2481 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.31+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_6' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='200*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='9.2e-07+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.089e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.4e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='4e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.85e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.31e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.7 nmos lmin=1.75e-07 lmax=1.85e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.608+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_7+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_7' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.57e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_7' ua='-2.032e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_7' ub='2.184e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_7' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_7' prwb=0.008 prwg=0.0 wr=1.0 u0='0.03416+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_7' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_7' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_7' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_7' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_7' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1943+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_7+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.548+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_7' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.5779 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1827 pdiblc1=0.1768 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03138 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.29+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_7' kt2=-0.02437 at=6.698e+4 ute=-1.53 ua1=6.012e-10 ub1=-3.37e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='200*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.189e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.2e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='3e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.78e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.01e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.15 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm02__model.8 nmos lmin=2.45e-07 lmax=2.55e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.599+sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_8+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_8' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.444e+05+sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_8' ua='-2.027e-09+sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_8' ub='2.272e-18+sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_8' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_8' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0299+sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_8' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_8' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_8' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_8' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_8' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.1943+sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_8+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='2.136+sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_8' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.5779 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1827 pdiblc1=0.1627 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.624e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03138 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.29+sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_8' kt2=-0.02437 at=6.698e+4 ute=-1.53 ua1=6.012e-10 ub1=-3.37e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='200*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.489e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='2e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='9e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.78e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.21e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.15 pbswgs=0.9064
.ends sky130_fd_pr__rf_nfet_01v8_bm02w5p00
.subckt sky130_fd_pr__rf_nfet_01v8_bm04 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_01v8_bm04 d g s b sky130_fd_pr__rf_nfet_01v8_bm04__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.0 nmos lmin=1.45e-07 lmax=1.55e-07 wmin=1.645e-06 wmax=1.655e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.90 rnoib=0.36 tnoia=2.7e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.604+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_0+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_0' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.744e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_0' ua='-1.96e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_0' ub='2.31e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_0' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_0' prwb=0.008 prwg=0.0 wr=1.0 u0='0.039+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_0' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_0' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_0' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_0' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_0' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.206+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_0+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='2.808+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_0' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.3121 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1748 pdiblc1=0.2729 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.29+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_0' kt2=-0.02437 at=5.978e+4 ute=-1.681 ua1=6.012e-10 ub1=-4.98e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='1800*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.083e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.559e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.64e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.58e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.91e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.1 nmos lmin=1.75e-07 lmax=1.85e-07 wmin=1.645e-06 wmax=1.655e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.90 rnoib=0.36 tnoia=2.7e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.6282+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_1+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_1' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_1' ua='-1.96e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_1' ub='2.31e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_1' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_1' prwb=0.008 prwg=0.0 wr=1.0 u0='0.036+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_1' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_1' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_1' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_1' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_1' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.206+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_1+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.685+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_1' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.3121 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1548 pdiblc1=0.1965 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03397 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.29+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_1' kt2=-0.02437 at=5.978e+4 ute=-1.681 ua1=6.012e-10 ub1=-4.98e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='1800*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.35e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.889e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.74e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.68e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.21e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.2 nmos lmin=2.45e-07 lmax=2.55e-07 wmin=1.645e-06 wmax=1.655e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.939e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.90 rnoib=0.36 tnoia=2.7e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=3.1e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.6095+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_2+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_2' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.544e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_2' ua='-2.02e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_2' ub='2.344e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_2' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_2' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0286+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_2' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_2' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_2' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_2' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_2' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.206+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_2+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='2.022+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_2' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.3121 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1548 pdiblc1=0.1965 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03397 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.29+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_2' kt2=-0.02437 at=5.978e+4 ute=-1.681 ua1=6.012e-10 ub1=-4.98e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='1800*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.35e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.989e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='4.04e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='8e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='1.0e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.68e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='1.81e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9064
.ends sky130_fd_pr__rf_nfet_01v8_bm04
.subckt sky130_fd_pr__rf_nfet_01v8_bm04w3p00 d g s b
.param l=1
.param w=3.01
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_01v8_bm04w3p00 d g s b sky130_fd_pr__rf_nfet_01v8_bm04__model l='l' w=3.01 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.3 nmos lmin=1.45e-07 lmax=1.55e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.076e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=2.2e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.593+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_3+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_3' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_3' ua='-2.032e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_3' ub='2.16e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_3' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_3' prwb=0.008 prwg=0.0 wr=1.0 u0='0.03499+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_3' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_3' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_3' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_3' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_3' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.2313+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_3+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='2.752+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_3' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.204 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1986 pdiblc1=0.19 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2112+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_3' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='880*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.274e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.069e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='3e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.7e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.21e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.4 nmos lmin=1.75e-07 lmax=1.85e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.076e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=2.2e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.612+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_4+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_4' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.594e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_4' ua='-2.032e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_4' ub='2.18e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_4' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_4' prwb=0.008 prwg=0.0 wr=1.0 u0='0.03129+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_4' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_4' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_4' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_4' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_4' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.2313+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_4+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.761+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_4' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.204 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1509 pdiblc1=0.1482 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2112+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_4' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='880*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.509e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.5e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.7e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='3.21e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.5 nmos lmin=2.45e-07 lmax=2.55e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.076e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=2.2e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.599+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_5+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_5' k3=3.0 dvt0=0.01 dvt1=0.2 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.498e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_5' ua='-2.052e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_5' ub='2.28e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_5' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_5' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0275+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_5' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_5' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_5' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_5' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_5' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.2313+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_5+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.902+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_5' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.204 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1177 pdiblc1=0.1363 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03202 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2112+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_5' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='880*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.809e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.8e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='7e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='9e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.7e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.21e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.ends sky130_fd_pr__rf_nfet_01v8_bm04w3p00
.subckt sky130_fd_pr__rf_nfet_01v8_bm04w5p00 d g s b
.param l=1
.param w=5.05
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_01v8_bm04w5p00 d g s b sky130_fd_pr__rf_nfet_01v8_bm04__model l='l' w=5.05 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.6 nmos lmin=1.45e-07 lmax=1.55e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.035e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=2.2e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.59+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_6+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_6' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.644e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_6' ua='-2.152e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_6' ub='2.44e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_6' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_6' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0354+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_6' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_6' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_6' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_6' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_6' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.2313+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_6+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='2.257+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_6' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.204 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1589 pdiblc1=0.1976 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03074 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2112+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_6' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='400*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.069e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='1e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.7e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.81e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.7 nmos lmin=1.75e-07 lmax=1.85e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.035e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=2.2e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.606+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_7+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_7' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.594e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_7' ua='-2.162e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_7' ub='2.461e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_7' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_7' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0314+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_7' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_7' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_7' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_7' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_7' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.2313+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_7+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.76+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_7' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.204 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1208 pdiblc1=0.1462 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03074 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2112+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_7' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='400*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.25e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.269e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.4e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='6e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.7e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.81e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.model sky130_fd_pr__rf_nfet_01v8_bm04__model.8 nmos lmin=2.45e-07 lmax=2.55e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.148e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='-2.035e-08+sky130_fd_pr__rf_nfet_01v8_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='9.181e-09+sky130_fd_pr__rf_nfet_01v8_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=0.0 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=-1.0e-7 vfbsdoff=0.0 lambda=0.0 vtl=2.0e+5 lc=5.0e-9 xn=3.0 rnoia=0.94 rnoib=0.26 tnoia=1.5e+7 tnoib=9.9e+6 epsrox=3.9 toxe='4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult+sky130_fd_pr__rf_nfet_01v8__b_toxe_slope_spectre*(4.148e-09*sky130_fd_pr__rf_nfet_01v8_b__toxe_mult*(sky130_fd_pr__rf_nfet_01v8__b_toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=2.2e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_01v8_b__rshg_diff' rsh=1.0 vth0='0.59+sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_8+sky130_fd_pr__rf_nfet_01v8__b_vth0_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_vth0_slope/sqrt(l*w*mult))' k1=0.5415 k2='-0.07197+sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_8' k3=3.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-0.2864 dvt1w=1.671e+6 dvt2w=-0.3571 w0=0.0 k3b=1.48 phin=0.0 lpe0=1.342e-7 lpeb=-7.224e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.524e+05+sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_8' ua='-2.102e-09+sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_8' ub='2.451e-18+sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_8' uc=7.917e-11 rdsw='98.95+sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_8' prwb=0.008 prwg=0.0 wr=1.0 u0='0.0274+sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_8' a0='1.471+sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_8' keta=0.1378 a1=0.0 a2=0.4239 ags='0.5074+sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_8' b0='-1.502e-07+sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_8' b1='1.902e-09+sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_8' eu=1.67 rdswmin=0.0 rdw=98.95 rdwmin=0.0 rsw=98.95 rswmin=0.0 voff='-0.2313+sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_8+sky130_fd_pr__rf_nfet_01v8__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_01v8__b_voff_slope/sqrt(l*w*mult))' nfactor='1.76+sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_8' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.204 etab=0.0001546 dsub=0.4657 voffl=5.82e-9 minv=0.0 pclm=0.1208 pdiblc1=0.1287 pdiblc2=0.0 pdiblcb=-1.0 drout=0.2457 pscbe1=3.295e+8 pscbe2=2.0e-6 pvag=0.0 delta=0.03074 alpha0=1.21e-7 alpha1=0.8767 beta0=14.77 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2.3e+9 cgidl=0.5 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=0.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.148e-9 kt1='-0.2112+sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_8' kt2=-0.02437 at=7.202e+4 ute=-1.681 ua1=6.012e-10 ub1=-7.32e-19 uc1=1.09e-12 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='400*sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult' rbpd=0.001 rbps=0.001 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.5e+42 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.84 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.3e-06+sky130_fd_pr__rf_nfet_01v8_b__xgw_diff' ngcon=2.0 diomod=1.0 njs=1.293 jss=0.00275 jsws=6.0e-10 xtis=2.0 bvs=11.9 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001229 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 cgdo='3.569e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgso='3.4e-10*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cgdl='8e-11*sky130_fd_pr__rf_nfet_01v8_b__overlap_mult' cf=1.0e-11 clc=1.2e-8 cle=1.9 dlc='2.3e-08+sky130_fd_pr__rf_nfet_01v8_b__dlc_diff+sky130_fd_pr__rf_nfet_01v8__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_01v8_b__dwc_diff' vfbcv=-1.0 acde=0.3801 moin=23.81 noff=1.0 voffcv=-0.06 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.0024*sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult' mjs=0.322 pbs=0.9877 cjsws='2.013e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjsws=0.001 pbsws=0.4 cjswgs='2.01e-10*sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult' mjswgs=0.1 pbswgs=0.9964
.ends sky130_fd_pr__rf_nfet_01v8_bm04w5p00