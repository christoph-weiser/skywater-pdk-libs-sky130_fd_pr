* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__slope=0.0
.subckt sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield c0 c1 b
.param mult=1.0
.param ctot_a='40.728e-15*sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor+1.06714/sqrt(mult/0.346925)*sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__slope*40.728e-15*sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor'
.param c0_sub='3.241e-15*cli2s_vpp'
.param c1_sub='1.307e-15*cli2s_vpp'
.param rat_m2=0.3761
.param rat_m1=0.3856
.param rat_li=0.2383
.param cap_m2='rat_m2*ctot_a'
.param cap_m1='rat_m1*ctot_a'
.param cap_li='rat_li*ctot_a'
.param lm2=3.685
.param wm2=0.140
.param nfm2=44.0
.param nvia_c0=84.0
.param nvia_c1=42.0
.param lm1=3.290
.param wm1=0.140
.param nfm1=52.0
.param ncon_c0=84.0
.param ncon_c1=16.0
.param ll1=3.655
.param wl1=0.170
.param nfl1=38.0
rm21 c0 a1 r='rm2*lm2/wm2*(1/3)*(1/nfm2)'
ccmvpp8p6x7p9 a1 c1 c='cap_m2'
rvia1 c0 d0 r='rcvia/nvia_c0'
rvia2 c1 d1 r='rcvia/nvia_c1'
rm11 d0 b1 r='rm1*lm1/wm1*(1/3)*(1/nfm1)'
cm1 b1 d1 c='cap_m1'
rcon1 d0 e0 r='rcl1/ncon_c0'
rcon2 d1 e1 r='rcl1/ncon_c1'
rli1 e0 f1 r='rl1*ll1/wl1*(1/3)*(1/nfl1)'
cli f1 e1 c='cap_li'
cli1_b e0 b c='c0_sub'
cli2_b e1 b c='c1_sub'
.ends sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield