* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8__toxe_slope=8.989e-03
.param sky130_fd_pr__rf_nfet_01v8__toxe1_slope=6.989e-03
.param sky130_fd_pr__rf_nfet_01v8__toxe2_slope=5.989e-03
.param sky130_fd_pr__rf_nfet_01v8__toxe3_slope=1.089e-02
.param sky130_fd_pr__rf_nfet_01v8__toxe4_slope=1.289e-02
.param sky130_fd_pr__rf_nfet_01v8__lint_slope=5.767e-9
.param sky130_fd_pr__rf_nfet_01v8__lint1_slope=0
.param sky130_fd_pr__rf_nfet_01v8__b_toxe_slope=3.443e-03
.param sky130_fd_pr__rf_nfet_01v8__b_voff_slope=0.007
.param sky130_fd_pr__rf_nfet_01v8__b_vth0_slope=5.556e-03