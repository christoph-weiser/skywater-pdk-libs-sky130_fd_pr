* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p84l0p15 d g s b
.param mult=1.0
.param rg_stub_tnom='(127*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult)'
.param rg_dist_tnom='(33.62*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p84l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(2)*(0.84)' ad='(2)*(0.1176)' as='(2)*(0.235)' pd='(2)*(1.12)' ps='(2)*(2.24)' nrd='(0)/(2)' nrs='(0)/(2)' nf=2 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(0.172f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gs 2 3 c='(0.07f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gd 2 1 c='(0.25f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(48*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(97*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p84l0p15
.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15 d g s b
.param mult=1.0
.param rg_stub_tnom='(63.5*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult)'
.param rg_dist_tnom='(16.81*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(4)*(0.84)' ad='(4)*(0.1176)' as='(4)*(0.176)' pd='(4)*(1.12)' ps='(4)*(1.68)' nrd='(0)/(4)' nrs='(0)/(4)' nf=4 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(0.41f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gs 2 3 c='(0.15f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gd 2 1 c='(0.59f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(32*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(50*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15
.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af04w3p00l0p15 d g s b
.param mult=1.0
.param rg_stub_tnom='(63.5*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult)'
.param rg_dist_tnom='(81.745*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af04w3p00l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(4)*(3.00)' ad='(4)*(0.42)' as='(4)*(0.63)' pd='(4)*(3.28)' ps='(4)*(4.92)' nrd='(0)/(4)' nrs='(0)/(4)' nf=4 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(1.47f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gs 2 3 c='(0.305f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gd 2 1 c='(0.73f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(8*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(14*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af04w3p00l0p15
.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15 d g s b
.param mult=1.0
.param rg_dist_nlrf_p42p15nf2=466.81
.param rg_stub_tnom='(127*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42)'
.param rg_dist_tnom='(rg_dist_nlrf_p42p15nf2*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(2)*(0.42)' ad='(2)*(0.0588)' as='(2)*(0.118)' pd='(2)*(0.7)' ps='(2)*(1.4)' nrd='(0)/(2)' nrs='(0)/(2)' nf=2 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(0.09f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42)'
cpar_gs 2 3 c='(0.115f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42)'
cpar_gd 2 3 c='(0.242f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(95.8*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(195*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af02w3p00l0p15 d g s b
.param mult=1.0
.param rg_stub_tnom='(127*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult)'
.param rg_dist_tnom='(191.46*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w3p00l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(2)*(3.00)' ad='(2)*(0.42)' as='(2)*(0.84)' pd='(2)*(3.28)' ps='(2)*(6.56)' nrd='(0)/(2)' nrs='(0)/(2)' nf=2 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(0.7f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gs 2 3 c='(0.163f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gd 2 1 c='(0.456f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(12*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(26*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af02w3p00l0p15
.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15 d g s b
.param mult=1.0
.param rg_stub_tnom='(31.75*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult)'
.param rg_dist_tnom='(40.87*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(8)*(3.00)' ad='(8)*(0.42)' as='(8)*(0.525)' pd='(8)*(3.28)' ps='(8)*(4.1)' nrd='(0)/(8)' nrs='(0)/(8)' nf=8 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(2.92f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gs 2 3 c='(0.61f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gd 2 1 c='(1.45f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(4.8*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(7*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15
.subckt sky130_fd_pr__rf_nfet_01v8_lvt_af08w0p84l0p15 d g s b
.param mult=1.0
.param rg_stub_tnom='(31.75*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult)'
.param rg_dist_tnom='(12.405*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult)'
.param tref=30.0
xsky130_fd_pr__rf_nfet_01v8_lvt_af08w0p84l0p15 1 2 3 b sky130_fd_pr__nfet_01v8_lvt l=0.15 w='(8)*(0.84)' ad='(8)*(0.1176)' as='(8)*(0.147)' pd='(8)*(1.12)' ps='(8)*(1.4)' nrd='(0)/(8)' nrs='(0)/(8)' nf=8 sa=0.28 sb=0.28 sd=0.28 m=1 mult='1*mult'
cpar_ds 1 3 c='(0.82f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gs 2 3 c='(0.33f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
cpar_gd 2 1 c='(0.84f*sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult)'
rg 2 g r='(rg_stub_tnom*(1+(temper-tref)*tc1rcgp+(temper-tref)*(temper-tref)*tc2rcgp))+(rg_dist_tnom*(1+(temper-tref)*tc1rsgpu+(temper-tref)*(temper-tref)*tc2rsgpu))'
rs 3 s r='(19.2*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult)'
rd 1 d r='(24.9*sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult)'
.ends sky130_fd_pr__rf_nfet_01v8_lvt_af08w0p84l0p15