* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_20v0__pwdrainjunction_mult=7.5058e-01
.param sky130_fd_pr__pfet_20v0__pwdrainmjswjunction_mult=8.3390e-1
.param sky130_fd_pr__pfet_20v0__pwdrainpbswjunction_mult=1.0204e+0
.param sky130_fd_pr__pfet_20v0__pwdrainctjunction_mult=1.0
.param sky130_fd_pr__pfet_20v0__vb=31.0
.param sky130_fd_pr__model__parasitic__diode_pw2dn__cj_mult=1.199716e+0
.param sky130_fd_pr__model__parasitic__diode_pw2dn__mj_mult=3.8681e-1
.param sky130_fd_pr__model__parasitic__diode_pw2dn__php_mult=1.0
.param sky130_fd_pr__model__parasitic__diode_pw2dn__tphp_mult=1.25
.param sky130_fd_pr__model__parasitic__diode_pw2dn__n_mult=1.0
.param sky130_fd_pr__model__parasitic__diode_pw2dn__js_mult=1.0
.model sky130_fd_pr__pfet_20v0__parasitic__diode_pw2dn d level=3.0 tlevc=1.0 scalm=1.0e-6 area=1.0e+12 cj='0.00038945*sky130_fd_pr__pfet_20v0__pwdrainjunction_mult*1e-12*sky130_fd_pr__model__parasitic__diode_pw2dn__ajunction_mult*sky130_fd_pr__model__parasitic__diode_pw2dn__cj_mult' mj='0.63982*sky130_fd_pr__pfet_20v0__pwdrainmjswjunction_mult*sky130_fd_pr__model__parasitic__diode_pw2dn__mj_mult' pb='0.58758*sky130_fd_pr__pfet_20v0__pwdrainpbswjunction_mult' cjsw='3.743e-010*sky130_fd_pr__pfet_20v0__pwdrainjunction_mult*1e-6*sky130_fd_pr__model__parasitic__diode_pw2dn__pjunction_mult*sky130_fd_pr__model__parasitic__diode_pw2dn__cj_mult' mjsw='0.80357*sky130_fd_pr__pfet_20v0__pwdrainmjswjunction_mult' php='0.2500*sky130_fd_pr__pfet_20v0__pwdrainpbswjunction_mult*sky130_fd_pr__model__parasitic__diode_pw2dn__php_mult' cta='0.0016157*sky130_fd_pr__pfet_20v0__pwdrainctjunction_mult' ctp='0.0008*sky130_fd_pr__pfet_20v0__pwdrainctjunction_mult' tpb=0.0010003 tphp='0.000675*sky130_fd_pr__model__parasitic__diode_pw2dn__tphp_mult' js='1.4693e-017*150' jsw='7.41e-018*150' n='1.0791*sky130_fd_pr__model__parasitic__diode_pw2dn__n_mult' rs=900 ik='2.08e-009/1e-12' ikr='0/1e-12' vb='sky130_fd_pr__pfet_20v0__vb' ibv=0.00106 trs=0 xti=3.0 eg=0.65 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0