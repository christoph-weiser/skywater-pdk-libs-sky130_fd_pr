* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_03v3_nvt__toxe_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__overlap_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__ajunction_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__pjunction_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__lint_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__wint_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__dlc_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__dwc_diff=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8=0.0
.include "sky130_fd_pr__nfet_03v3_nvt.pm3.spice"