* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_hvt__toxe_mult=0.9635
.param sky130_fd_pr__pfet_01v8_hvt__rshp_mult=1.0
.param sky130_fd_pr__pfet_01v8_hvt__overlap_mult=0.91216
.param sky130_fd_pr__pfet_01v8_hvt__lint_diff=1.21275e-8
.param sky130_fd_pr__pfet_01v8_hvt__wint_diff=-2.252e-8
.param sky130_fd_pr__pfet_01v8_hvt__dlc_diff=1.21275e-8
.param sky130_fd_pr__pfet_01v8_hvt__dwc_diff=-2.252e-8
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_0=1.1685
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_0=-0.073198
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_0=-0.0026118
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_0=9.5527e-20
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_0=0.00050729
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_0=-19944.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_0=-0.0030954
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_0=4.0273e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_0=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_1=1.3432
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_1=-0.092546
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_1=-1.9333e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_1=-0.012028
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_1=0.00091138
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_1=-9676.4
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_1=-0.031374
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_1=3.0168e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_2=0.56345
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_2=-0.10583
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_2=0.14627
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_2=-0.045106
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_2=3.3308e-21
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_2=-0.0032344
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_2=0.0017886
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_2=0.019608
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_2=2.0826e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_3=-4.0534e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_3=0.38734
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_3=-0.065774
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_3=0.07242
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_3=-0.033589
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_3=3.0272e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_3=-0.0065218
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_3=0.0015153
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_3=0.02967
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_3=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_4=-4.1332e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_4=0.31876
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_4=-0.055948
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_4=0.12352
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_4=-0.051614
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_4=2.6481e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_4=-0.0085758
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_4=0.0012323
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_4=0.023235
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_4=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_5=1.3844e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_5=0.42843
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_5=-0.016079
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_5=0.017163
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_5=-0.053143
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_5=2.3908e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_5=-0.0095913
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_5=0.0015095
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_5=0.021084
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_6=5.2669e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_6=1.9958
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_6=-0.12259
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_6=-3.4027e-19
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_6=-0.019713
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_6=0.0018756
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_6=-15042.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_6=-0.032438
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_7=0.00049592
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_7=3.6023e-19
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_7=10368.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_7=-0.042677
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_7=-1.069e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_7=0.67102
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_7=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_7=-0.088953
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_7=0.00628
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_8=0.0031239
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_8=0.0010265
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_8=2.1389e-19
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_8=-12024.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_8=0.027597
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_8=1.7824e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_8=0.7444
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_8=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_8=-0.041554
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_9=-0.064005
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_9=-0.011158
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_9=0.0033537
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_9=-9.374e-20
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_9=-1068.6
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_9=0.035019
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_9=5.9079e-10
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_9=0.81734
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_10=5.4485e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_10=-0.062192
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_10=0.030386
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_10=-0.077196
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_10=0.067058
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_10=0.0017933
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_10=0.014942
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_10=-0.01012
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_10=-1.423e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_11=-1.8151e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_11=7.7975e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_11=-0.059985
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_11=0.0073573
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_11=-0.017776
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_11=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_11=0.19926
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_11=0.0027314
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_11=0.012664
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_11=-0.010653
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_12=-0.01065
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_12=-1.2211e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_12=8.7918e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_12=-0.058568
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_12=0.11377
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_12=-0.073942
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_12=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_12=0.22168
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_12=0.0037612
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_12=-0.020239
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_13=0.17176
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_13=0.0040371
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_13=-0.00070285
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_13=-0.0082896
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_13=-2.9883e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_13=1.1918e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_13=-0.059659
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_13=0.082174
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_13=-0.048602
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_13=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_14=-14280.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_14=0.84074
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_14=0.00022368
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_14=-0.016864
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_14=-0.0070323
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_14=1.3205e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_14=5.1491e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_14=-0.095817
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_14=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_15=15711.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_15=0.65106
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_15=0.0012414
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_15=-0.049467
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_15=-0.0066346
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_15=2.433e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_15=-1.3804e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_15=-0.075268
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_15=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_16=-18555.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_16=0.80575
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_16=0.0015763
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_16=-0.0047728
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_16=0.0014215
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_16=2.4851e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_16=5.9683e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_16=-0.032169
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_16=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_17=0.29713
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_17=0.0021483
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_17=36492.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_17=0.012625
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_17=-0.0068541
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_17=8.7197e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_17=3.6509e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_17=-0.062892
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_17=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_18=0.042277
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_18=-0.054963
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_18=0.096808
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_18=0.0018384
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_18=0.011981
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_18=-0.011668
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_18=-1.3486e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_18=5.6391e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_18=-0.0579
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_19=-0.06713
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_19=0.089035
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_19=-0.09226
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_19=0.07946
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_19=0.0025237
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_19=-8.9723e-5
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_19=-0.0081353
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_19=-2.336e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_19=8.0784e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_20=-0.060164
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_20=0.05552
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_20=-0.060337
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_20=0.13939
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_20=0.0038347
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_20=-0.0013833
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_20=-0.0075985
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_20=-2.8979e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_20=1.1254e-18
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_21=1.0194e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_21=-0.040412
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_21=0.031765
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_21=-0.016859
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_21=0.16995
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_21=0.0035046
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_21=0.014807
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_21=-0.0064282
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_21=-2.7503e-10
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_22=2.8009e-12
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_22=1.0413e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_22=-0.061149
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_22=-16814.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_22=0.726
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_22=8.9971e-5
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_22=-0.036158
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_22=-0.003578
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_23=0.00078982
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_23=3.2854e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_23=-1.1949e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_23=-0.031663
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_23=-1225.1
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_23=0.77276
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_23=0.001374
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_23=-0.029264
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_24=0.19194
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_24=0.00055265
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_24=-0.0071206
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_24=2.4031e-5
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_24=-5.5968e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_24=2.8948e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_24=-0.042475
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_24=937.61
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_25=17793.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_25=0.035627
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_25=-3.0258e-5
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_25=0.024752
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_25=-0.0083859
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_25=-4.7515e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_25=8.3215e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_25=-0.047352
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_25=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_26=-0.057758
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_26=0.0028982
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_26=0.0026436
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_26=-0.0095685
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_26=-2.3523e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_26=8.6273e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_26=-0.061638
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_26=0.070775
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_26=-0.090391
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_26=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_27=-0.042836
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_27=0.0038855
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_27=0.00012138
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_27=-0.009744
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_27=-3.1095e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_27=1.1464e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_27=-0.049907
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_27=0.093034
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_27=-0.1001
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_27=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_28=0.13257
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_28=0.0038659
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_28=0.01494
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_28=-0.006178
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_28=-3.3863e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_28=1.1922e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_28=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_28=-0.042942
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_28=0.038848
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_28=-0.018152
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_29=0.031036
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_29=-0.022185
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_29=0.12009
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_29=0.0045545
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_29=0.0086119
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_29=-0.0097198
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_29=-3.5005e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_29=1.3167e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_29=-0.044302
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_30=-0.061481
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_30=-7933.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_30=1.0735
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_30=0.0013729
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_30=-0.045176
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_30=-0.025226
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_30=4.3641e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_30=-3.5991e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_31=-0.06935
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_31=10246.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_31=0.29389
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_31=-7.5611e-6
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_31=-0.058017
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_31=-0.0026065
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_31=-1.2333e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_31=2.3325e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_32=1.962e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_32=-0.054434
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_32=969.47
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_32=0.23975
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_32=0.00037356
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_32=-0.0015635
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_32=-0.00068126
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_32=-2.7637e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_33=1.9454e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_33=4.0906e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_33=-0.038333
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_33=-24495.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_33=0.77191
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_33=0.0018039
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_33=0.0099204
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_33=-0.0093591
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_34=-0.010952
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_34=2.3169e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_34=9.8491e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_34=-0.10242
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_34=-1.07e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_34=3.7245e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_34=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_34=1.1946
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_34=0.0065629
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_34=0.024445
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_35=0.33573
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_35=0.0030529
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_35=-0.018917
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_35=-0.014777
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_35=-2.1406e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_35=8.0918e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_35=-0.082328
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_35=-1.2969e-7
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_35=5.9733e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_36=0.46808
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_36=0.0041521
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_36=-0.00080103
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_36=-0.014506
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_36=-1.831e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_36=1.0548e-18
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_36=-0.088243
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_36=-2.3704e-9
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_36=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_36=3.9067e-10
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_37=3.1021e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_37=0.38657
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_37=0.0016757
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_37=0.024333
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_37=-0.0082481
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_37=-1.2102e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_37=3.7977e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_37=-0.064468
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_37=4.9916e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_37=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_38=9.7817e-9
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_38=-1.0548e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_38=0.33142
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_38=0.0018676
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_38=-0.00065254
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_38=-0.01054
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_38=-9.1285e-11
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_38=3.4787e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_38=-0.068041
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_38=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_39=1.5108
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_39=0.0014121
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_39=-33268.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_39=0.049605
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_39=-0.0033833
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_39=1.9943e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_39=2.4461e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_39=-0.17534
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_39=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_40=-20502.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_40=1.2981
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_40=0.0011093
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_40=0.013628
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_40=-0.011097
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_40=1.589e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_40=1.4831e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_40=-0.16376
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_40=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_41=-0.080356
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_41=-22215.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_41=1.2353
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_41=0.0048634
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_41=0.072171
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_41=-0.020607
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_41=3.7921e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_41=5.3941e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_42=-0.079199
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_42=3.312e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_42=-3.5189e-9
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_42=0.84927
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_42=0.0038212
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_42=0.022241
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_42=-0.013114
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_42=5.9893e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_42=-1.5614e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_43=2.4113e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_43=-0.052516
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_43=5.6987e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_43=6.3971e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_43=0.4197
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_43=0.0016695
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_43=0.0331
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_43=-0.0038093
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_43=2.2378e-11
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_44=-4.704e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_44=3.6014e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_44=-0.057818
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_44=3.7587e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_44=-9.6801e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_44=0.38267
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_44=0.0019947
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_44=0.023572
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_44=-0.0061834
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_45=-0.00737
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_45=-1.6303e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_45=4.1509e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_45=-0.054064
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_45=2.8315e-8
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_45=8.6241e-10
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_45=0.28425
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_45=0.0014955
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_45=0.018605
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_46=1.6519
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_46=0.0015386
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_46=-0.027131
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_46=-0.022499
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_46=3.2587e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_46=-5.8085e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_46=-0.10259
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_46=-27255.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_47=-46144.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_47=1.8927
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_47=0.0047167
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_47=0.065178
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_47=-0.0040734
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_47=2.546e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_47=8.0887e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_47=-0.069708
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_47=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_48=-10711.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_48=1.8855
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_48=0.00050012
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_48=-0.00043113
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_48=-0.0078901
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_48=-5.7141e-12
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_48=2.338e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_48=-0.16453
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_48=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_49=-15166.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_49=1.7817
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_49=0.0026371
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_49=0.0046864
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_49=-0.013314
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_49=8.0263e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_49=-4.6705e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_49=-0.11746
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_49=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_50=-16132.59856887
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_50=0.00053206
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_50=1.07943065
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_50=-0.01847513
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_50=0.00052558
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_50=8.10068e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_50=7.43303e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_50=-0.07226901
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_50=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_51=-4026.02605404
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_51=-0.00016362
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_51=0.55331993
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_51=-0.04239203
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_51=0.00420768
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_51=-2.4623e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_51=-1.9168e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_51=-0.054493
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_51=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_52=-0.04175202
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_52=-13981.97902176
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_52=0.0006674
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_52=0.8647004
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_52=-0.03223565
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_52=0.00575
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_52=1.7979e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_52=-9.8029e-20
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_52=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_53=-0.06030202
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_53=-2249.59441703
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_53=-0.00015602
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_53=0.73462969
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_53=-0.04329494
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_53=0.00426399
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_53=-4.418e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_53=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_53=3.569e-20
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_54=-5.4309e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_54=-0.068457
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_54=-9019.51550916
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_54=0.00244428
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_54=0.36719917
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_54=-0.04347459
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_54=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_54=-0.003124
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_54=8.10566e-10
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_55=2.57865e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_55=-2.21824e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_55=-0.017588
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_55=-17212.99898427
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_55=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_55=0.00070886
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_55=0.52491998
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_55=-0.04055681
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_55=0.0067584
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_56=-0.012919
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_56=5500.8
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_56=-0.00052794
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_56=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_56=0.067192
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_57=-0.00020347
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_57=0.010711
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_57=-0.0029141
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_57=-16610.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_57=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_58=-14143.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_58=-0.00024178
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_58=0.0047006
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_58=-0.0041664
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_58=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_59=-10943.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_59=0.00103419
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_59=0.001143
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_59=0.82063676
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_59=-0.026214
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_59=-0.011373
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_59=3.41926e-10
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_59=-1.46571e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_59=-0.00019276
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_59=-0.00097934
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_59=-0.07107368
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_59=3.08149e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_59=-5.0961e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_59=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_60=-5.23507e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_60=-7871.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_60=0.0015088
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_60=0.00106239
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_60=0.63824361
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_60=-0.032868
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_60=-0.011761
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_60=5.28643e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_60=-3.04591e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_60=-0.00019801
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_60=-0.07010265
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_60=-0.00100604
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_60=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_60=3.16552e-12
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_61=2.16233e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_61=-3.57602e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_61=-5364.7
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_61=0.00072571
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_61=0.0018234
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_61=0.50977511
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_61=-0.036338
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_61=-0.012049
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_61=6.61595e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_61=-4.17079e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_61=-0.00013526
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_61=-0.06935327
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_61=-0.00068722
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_61=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_62=9.63646e-13
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_62=-1.59366e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_62=-3473.1
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_62=0.00032341
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_62=0.0020537
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_62=0.42204309
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_62=-0.037835
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_62=-0.010776
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_62=7.53084e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_62=-4.94471e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_62=-6.02786e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_62=-0.06880988
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_62=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_62=-0.00030626
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_63=-0.00030626
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_63=-0.06880988
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_63=9.63645e-13
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_63=-1.59368e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_63=-5939.8
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_63=0.00032341
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_63=0.002182
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_63=0.42204238
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_63=-0.024116
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_63=-0.017273
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_63=7.53084e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_63=-4.94471e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_63=-6.02787e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_63=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_64=-8.28307e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_64=-311277.85910916
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_64=-0.00033188
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_64=0.00033957
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_64=-0.01854726
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_64=1.11822e-12
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_64=2.48144e-5
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_64=1733.5
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_64=0.0011099
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_64=0.24978359
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_64=0.015004
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_64=0.0015805
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_64=2.17866e-11
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_64=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_64=2.72104e-19
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_65=18392.0
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_65=-0.00019188
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_65=0.033219
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_65=-0.0034405
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_65=0.0
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_66=7.18929e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_66=-4.78344e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_66=0.00022885
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_66=-0.0645413
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_66=-3.24613e-13
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_66=1.37064e-6
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_66=2082.7
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_66=0.0
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_66=0.0019666
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_66=0.44034087
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_66=-0.039363
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_66=-0.010451
.param sky130_fd_pr__pfet_01v8_hvt__k2_diff_67=-0.0083591
.param sky130_fd_pr__pfet_01v8_hvt__rdsw_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__pdits_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ua_diff_67=3.91251e-10
.param sky130_fd_pr__pfet_01v8_hvt__pclm_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ub_diff_67=-2.47071e-19
.param sky130_fd_pr__pfet_01v8_hvt__kt1_diff_67=5.69173e-5
.param sky130_fd_pr__pfet_01v8_hvt__bgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__tvoff_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__cgidl_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__ags_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__a0_diff_67=0.00041074
.param sky130_fd_pr__pfet_01v8_hvt__voff_diff_67=-0.05063977
.param sky130_fd_pr__pfet_01v8_hvt__pditsd_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__agidl_diff_67=-5.82603e-13
.param sky130_fd_pr__pfet_01v8_hvt__keta_diff_67=2.46002e-6
.param sky130_fd_pr__pfet_01v8_hvt__b0_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__b1_diff_67=0.0
.param sky130_fd_pr__pfet_01v8_hvt__vsat_diff_67=3559.7
.param sky130_fd_pr__pfet_01v8_hvt__eta0_diff_67=3.3371e-5
.param sky130_fd_pr__pfet_01v8_hvt__u0_diff_67=0.0010084
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_diff_67=0.6994729
.param sky130_fd_pr__pfet_01v8_hvt__vth0_diff_67=-0.028431
.include "sky130_fd_pr__pfet_01v8_hvt__ff.pm3.spice"