* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8_lvt__toxe_mult=0.9635
.param sky130_fd_pr__nfet_01v8_lvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8_lvt__overlap_mult=0.88119
.param sky130_fd_pr__nfet_01v8_lvt__ajunction_mult=0.87784
.param sky130_fd_pr__nfet_01v8_lvt__pjunction_mult=0.78244
.param sky130_fd_pr__nfet_01v8_lvt__lint_diff=1.21275e-8
.param sky130_fd_pr__nfet_01v8_lvt__wint_diff=-2.252e-8
.param sky130_fd_pr__nfet_01v8_lvt__dlc_diff=7.7131e-9
.param sky130_fd_pr__nfet_01v8_lvt__dwc_diff=-2.252e-8
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_0=-0.064001
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_0=0.0081134
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_0=0.0020103
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_0=-0.10975
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_0=-7.0587e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_0=3.8853e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0=0.70456
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0=-0.0076786
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_1=-0.050662
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_1=0.0077884
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_1=-0.10908
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_1=0.00093901
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_1=6.8072e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_1=2.826e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1=0.39852
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1=-0.0078928
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2=-0.0043298
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_2=0.0090734
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_2=0.0099409
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_2=-0.0061366
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_2=0.00062214
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_2=-1.9272e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_2=2.575e-19
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2=0.72829
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3=1.4729
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3=-0.058087
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_3=0.031103
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_3=-0.0015859
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_3=6.8273e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3=-26072.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_3=1.612e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4=1.5178
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4=-0.082199
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_4=0.019857
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_4=-0.0021861
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_4=1.8015e-11
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4=-21912.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_4=4.5553e-20
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_5=4.5063e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5=0.95603
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5=-0.011184
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_5=0.0093294
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_5=0.0024348
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_5=-2.0398e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5=-12947.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_6=2.7444e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6=1.3429
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6=-0.010655
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_6=-0.00062272
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_6=0.0005695
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_6=-3.92e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6=-10142.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_7=2.4261e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7=0.77503
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7=8.7015e-5
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_7=-0.026006
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_7=0.0038481
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_7=-0.035935
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_7=0.0013497
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_7=-2.3833e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_8=-0.034253
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_8=0.00070921
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_8=-5.0806e-13
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_8=1.9943e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8=0.36129
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8=-0.0057838
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_8=-0.020934
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_8=0.0013629
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_9=-0.006192
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_9=0.00026333
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_9=-1.1842e-12
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_9=1.3971e-19
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9=0.42662
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9=-0.00025391
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_9=0.0058881
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_9=0.0058275
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_10=3.5409e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_10=-1.1456e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_10=-0.0028995
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10=-19021.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10=-0.085201
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10=1.2225
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_10=0.033776
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_11=0.024793
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_11=2.1273e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_11=1.6509e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_11=-0.00039822
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11=-12938.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11=-0.063158
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11=1.2006
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_12=0.014212
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_12=-8.5273e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_12=4.9607e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_12=0.0012429
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12=-7928.4
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12=-0.020197
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12=0.93234
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_13=0.012015
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_13=9.2164e-14
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_13=2.3157e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_13=0.00020896
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13=-6126.5
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13=-0.0076636
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13=1.2266
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14=0.63062
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_14=0.0029183
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_14=-1.0862e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_14=2.207e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_14=-0.033478
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_14=-0.050039
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_14=0.00097848
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14=-0.0082701
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15=0.00092243
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15=0.51633
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_15=-0.0060606
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_15=-1.8742e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_15=2.3666e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_15=0.011196
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_15=0.015378
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_15=0.00093567
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_16=-0.02206
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_16=0.00051071
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16=-0.010136
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16=0.10272
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_16=0.0085836
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_16=1.3225e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_16=1.6378e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_16=0.0031853
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_17=-0.00082717
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17=-13818.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17=-0.074175
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17=1.3395
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_17=0.037049
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_17=2.9203e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_17=1.1213e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_18=-0.0012159
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18=-16297.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18=-0.047066
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18=1.2712
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_18=0.025327
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_18=2.6552e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_18=8.029e-20
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_19=3.6615e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_19=0.00042198
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19=-13450.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19=-0.028005
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19=0.75655
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_19=0.011293
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_19=-3.8741e-11
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_20=-2.0719e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_20=2.5573e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_20=0.00081091
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20=-899.91
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20=-0.011093
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20=1.1478
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_20=0.0019437
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_21=-4.2056e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_21=2.5388e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_21=0.045409
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_21=0.048057
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_21=0.0013807
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21=0.00038533
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21=0.74534
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_21=-0.0047384
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_22=0.0076765
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_22=-1.281e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_22=1.9584e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_22=0.00072066
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_22=-0.0067956
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_22=0.00074354
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22=-0.0053605
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22=0.45602
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_23=0.0067583
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_23=-2.3598e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_23=2.1315e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_23=-0.00059699
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_23=0.031865
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_23=0.0010023
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23=-0.004118
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23=0.3288
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_24=0.038683
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_24=1.1967e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_24=-1.6049e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_24=-0.0047096
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24=-14167.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24=-0.089849
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24=1.3376
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25=1.2419
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_25=0.022825
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_25=6.4936e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_25=-2.5046e-21
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_25=-0.0023153
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25=-15924.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25=-0.046521
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26=-0.018801
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26=0.73783
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_26=0.01227
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_26=-1.2398e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_26=3.5666e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_26=0.0014372
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26=-11322.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_27=0.00066763
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27=-1962.1
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27=-0.0048024
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27=0.98774
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_27=0.0037101
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_27=-2.8272e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_27=2.1671e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_28=0.002882
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28=-0.018416
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28=0.13245
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_28=9.6413e-8
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_28=1.0459e-9
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_28=0.0046606
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_28=-1.7631e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_28=5.0687e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_29=-0.0019238
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29=-26661.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29=-0.11716
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29=1.6054
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_29=0.029703
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_29=4.346e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_29=1.5069e-19
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_30=6.8804e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_30=-0.00058909
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30=-22958.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30=-0.10542
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30=1.5302
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_30=0.012433
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_30=2.2286e-11
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_31=2.689e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_31=-3.4876e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_31=-0.0029007
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31=-34751.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31=-0.13397
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31=2.1416
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_31=0.017083
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_32=2.0615e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_32=3.0798e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_32=-0.0015571
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32=-19624.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32=-0.13512
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32=2.159
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_32=0.017306
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_33=0.016181
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_33=2.0951e-11
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_33=-7.6709e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_33=-0.0019419
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33=-15572.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33=-0.12569
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33=1.9124
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_34=0.031783
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_34=1.2373e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_34=-1.044e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_34=-0.0033755
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34=-17260.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34=-0.087483
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34=1.646
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_35=0.032894
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_35=2.3003e-12
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_35=-7.6801e-20
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_35=-0.0030264
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35=-21178.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35=-0.083109
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35=1.2691
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36=1.4374
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_36=0.037302
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_36=9.319e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_36=1.7106e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_36=-0.00099139
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36=-13868.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36=-0.071658
.param sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37=-0.023221
.param sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37=0.89187
.param sky130_fd_pr__nfet_01v8_lvt__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__b1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__k2_diff_37=0.010877
.param sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ua_diff_37=-2.1819e-13
.param sky130_fd_pr__nfet_01v8_lvt__ub_diff_37=3.2503e-19
.param sky130_fd_pr__nfet_01v8_lvt__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8_lvt__u0_diff_37=0.00072118
.param sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37=-12287.0
.include "sky130_fd_pr__nfet_01v8_lvt.pm3.spice"