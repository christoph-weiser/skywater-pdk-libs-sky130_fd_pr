* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param tol_nfom=0.069u
.param tol_pfom=0.060u
.param tol_nw=0.069u
.param tol_poly=0.041u
.param tol_li=0.020u
.param tol_m1=0.025u
.param tol_m2=0.025u
.param tol_m3=0.065u
.param tol_m4=0.065u
.param tol_m5=0.17u
.param tol_rdl=1.0u
.param rcn=70
.param rcp=330
.param rdn=108
.param rdp=166
.param rdn_hv=102
.param rdp_hv=160
.param rp1=42.2
.param rnw=1240
.param rl1=9.5
.param rm1=0.105
.param rm2=0.105
.param rm3=0.038
.param rm4=0.038
.param rm5=0.0212
.param rrdl=0.004
.param rcp1=25.28
.param rcl1=1.6
.param rcvia=2.0
.param rcvia2=0.50
.param rcvia3=0.50
.param rcvia4=0.012
.param rcrdlcon=0.0046
.param rspwres=2803
.param crpf_precision=1.53e-04
.param crpfsw_precision_1_1=5.83e-11
.param crpfsw_precision_2_1=6.19e-11
.param crpfsw_precision_4_1=6.66e-11
.param crpfsw_precision_8_2=7.22e-11
.param crpfsw_precision_16_2=7.88e-11
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/slow.spice"