* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__cap_var_lvt c0 c1 b w=5 l=0.5 vm=1 wc='w*1' lc='l*1'
.param cnwvc_ldiff=0.15
.param wd='wc+2*cnwvc_dwc'
.param ld='lc+2*cnwvc_dlc'
.param ldd='0.018+2*cnwvc_dld'
.param dwr=-0.02
.param dwp=-0.5
.param dlr=0.02
.param wl='(wd-2*dwr)/(ld-2*dlr)'
.param wlwdiff='((0.5*(ld-2*dlr))+cnwvc_ldiff)/(2*(wd-2*dwr))'
.param sky130_fd_pr__cap_var_lvt__cmin_slope_l=1.1e-16
.param sky130_fd_pr__cap_var_lvt__cmin_slope_w=1.5e-16
.param sky130_fd_pr__cap_var_lvt__cmin_slope_wl=3.5e-16
.param sky130_fd_pr__cap_var_lvt__cmax_slope_l=7.0e-16
.param sky130_fd_pr__cap_var_lvt__cmax_slope_w=7.0e-16
.param sky130_fd_pr__cap_var_lvt__cmax_slope_wl=1.5e-15
.param cnwvc_slope1=0.21875
.param cnwvc_slope2=0.125
.param cm0='5.571e-16*cnwvc_cintmult'
.param cm1='4.775e-16'
.param dev/gauss='sky130_fd_pr__cap_var_lvt__cmin_slope_l/sqrt(2*ld*vm)'
.param cm2='2.019e-16'
.param dev/gauss='sky130_fd_pr__cap_var_lvt__cmin_slope_w/sqrt(2*wd*vm)'
.param cm3='6.529e-16*cnwvc_cdepmult'
.param dev/gauss='sky130_fd_pr__cap_var_lvt__cmin_slope_wl*cnwvc_cdepmult/sqrt(2*ld*wd*vm)'
.param cx0=6.261e-16
.param cx1='5.75e-16'
.param dev/gauss='sky130_fd_pr__cap_var_lvt__cmax_slope_l/sqrt(2*ld*vm)'
.param cx2='1.712e-16'
.param dev/gauss='sky130_fd_pr__cap_var_lvt__cmax_slope_w/sqrt(2*wd*vm)'
.param cx3='8.854e-14*3.9/cnwvc_tox'
.param dev/gauss='sky130_fd_pr__cap_var_lvt__cmax_slope_wl/sqrt(2*wd*ld*vm)'
.param sky130_fd_pr__cap_var_lvt__vgs_min_1='-2.071'
.param sky130_fd_pr__cap_var_lvt__vgs_max_1='-1*-2.071'
.param sky130_fd_pr__cap_var_lvt__tmax_vgs_1='100.001n'
.param sky130_fd_pr__cap_var_lvt__vgs_min_2='-2.161'
.param sky130_fd_pr__cap_var_lvt__vgs_max_2='-1*-2.161'
.param sky130_fd_pr__cap_var_lvt__tmax_vgs_2='20.001n'
.param sky130_fd_pr__cap_var_lvt__vgs_min='-2.301'
.param sky130_fd_pr__cap_var_lvt__vgs_max='-1*-2.301'
.param tref=30.0
.param cmin='cm0+cm1*ld+cm2*wd+cm3*wd*(ld-ldd)+cx3*wd*ldd'
.param cmax='cx0+cx1*ld+cx2*wd+cx3*wd*ld'
cg c0 p2 q='cmin*vm*(v(c0)-v(p2))+((0.5*(cmax+cmin)-cmin)*(v(c0)-v(p2))+0.5*(cmax-cmin)*(1/1.9)*(cnwvc_slope1*log(cosh((v(c0)-v(p2)-cnwvc_vt1)/cnwvc_slope1))+0.9*cnwvc_slope2*log(cosh((v(c0)-v(p2)-cnwvc_vt2)/cnwvc_slope2))))*vm'
c3 c0 b c='0.15e-15'
c4 c1 b c='0.15e-15'
.param con_sp=0.17
.param cnwvc_k=12
.param cnwvc_n1=0.1
.param cnwvc_n2=0.28
.param apoly=1.15
.param apolyc=1
.param acon=1
.param anwell=1
.param bnwell=0.6
.param cnwell=2
.param n_pocon='max((lc-0.14)/(2*con_sp),1)'
.param n_con='(wc-2*0.06+con_sp)/(2*con_sp)'
.param rg_tc1=3e-3
.param rg_tc2=0.0
.param rg_tcmult='1+(temper-tref)*rg_tc1+(temper-tref)*(temper-tref)*rg_tc2'
.param cnwvc_a='apoly*rp1*wl/cnwvc_k+apolyc*rcp1/n_pocon+acon*rcn/n_con+anwell*rnw*wlwdiff'
.param cnwvc_b1='bnwell*rnw*wlwdiff'
.param cnwvc_c='cnwell*rnw*((0.5*(ld-2*dlr))+cnwvc_ldiff)/(2*(wd-2*dwp))'
rg p2 c1 r='(cnwvc_a+cnwvc_b1*(0.5*tanh((v(c0)-v(p2)-cnwvc_vtr)/cnwvc_n1)+0.5)+20*cnwvc_c*(0.5*tanh((v(c0)-v(p2)-cnwvc_vtr)/cnwvc_n1)+0.5)*exp(-abs((v(c0)-v(p2)-cnwvc_vtr)/cnwvc_n2)))/vm*rg_tcmult'
.ends sky130_fd_pr__cap_var_lvt