* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_g5v0d10v5__toxe_mult=0.94
.param sky130_fd_pr__nfet_g5v0d10v5__rshn_mult=1.0
.param sky130_fd_pr__nfet_g5v0d10v5__overlap_mult=0.76246
.param sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult=0.81753
.param sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult=0.77786
.param sky130_fd_pr__nfet_g5v0d10v5__lint_diff=1.7325e-8
.param sky130_fd_pr__nfet_g5v0d10v5__wint_diff=-3.2175e-8
.param sky130_fd_pr__nfet_g5v0d10v5__dlc_diff=1.7325e-8
.param sky130_fd_pr__nfet_g5v0d10v5__dwc_diff=-3.2175e-8
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_0=-0.001744
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_0=0.00067346
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_0=-0.11661
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_0=-0.18148
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_0=-7.2729e-13
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_0=-10837.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_0=-0.31653
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_0=-8.9194e-20
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_1=0.0065028
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_1=-0.00072595
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_1=-0.038431
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_1=-2.7173e-11
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_1=-0.17178
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_1=-0.36457
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_1=-2.9245e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_1=0.096329
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_1=-0.27221
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_1=-5.5898e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_2=-0.33559
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_2=-2.1053e-19
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_2=-0.0025359
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_2=0.0018816
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_2=-0.10427
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_2=3.0e-7
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_2=-0.20323
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_2=-6.098e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_2=-6890.7
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_3=0.24311
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_3=-2.8366e-19
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_3=-0.0024725
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_3=-0.0031377
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_3=-0.06814
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_3=1.7281e-6
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_3=-0.11561
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_3=-0.09111
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_3=3.524e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_3=0.041256
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_4=0.0010053
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_4=0.53181
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_4=-2.4973e-19
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_4=-0.012359
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_4=-0.0025723
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_4=-0.042806
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_4=3.1541e-11
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_4=-0.019831
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_4=-0.15691
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_4=2.6852e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_5=2.0835e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_5=0.0022408
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_5=-1.6048e-19
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_5=0.57949
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_5=-0.015725
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_5=-0.0016407
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_5=-0.023815
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_5=1.2456e-10
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_5=-0.018345
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_5=-0.37378
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_6=-0.13163
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_6=9.6095e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_6=-17518.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_6=2.1831e-19
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_6=-0.17311
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_6=0.0086273
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_6=-0.0017875
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_6=-0.15352
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_6=3.0e-7
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_7=6.9949e-7
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_7=-0.53824
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_7=-0.080439
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_7=9.0617e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_7=-0.59992
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_7=-4.0753e-20
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_7=0.30855
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_7=0.005737
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_7=-0.00061823
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_7=-0.051511
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_8=-0.045086
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_8=-0.19936
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_8=2.8087e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_8=0.0065931
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_8=3.9997e-20
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_8=0.55919
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_8=-0.01817
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_8=-0.00080585
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_8=-0.040256
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_8=6.5034e-11
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_9=1.8224e-10
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_9=-0.0012822
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_9=-0.05098
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_9=-0.42307
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_9=1.4474e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_9=0.0068253
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_9=-1.5723e-19
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_9=0.59935
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_9=-0.011513
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_9=-0.029635
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_10=0.0033427
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_10=-0.00063338
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_10=-0.020704
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_10=1.8393e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_10=-0.02635
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_10=-0.013333
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_10=-0.56346
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_10=0.94736
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_10=1.0675e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_10=3.155e-20
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_11=-0.11536
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_11=6.1171e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_11=-0.0015314
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_11=-16625.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_11=-0.13341
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_11=0.012032
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_11=-0.10634
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_11=1.6344e-11
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_12=-0.12
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_12=5.7445e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_12=-0.16844
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_12=2.1575e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_12=-0.00080036
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_12=-16866.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_12=3.8187e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_12=-0.099541
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_12=0.00028865
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_13=-0.0036231
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_13=0.015715
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_13=5.462e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_13=-0.27985
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_13=1.5753e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_13=-0.0011108
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_13=-15059.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_13=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_13=2.9615e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_13=-0.051577
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_14=-0.033955
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_14=0.0059175
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_14=-0.042183
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_14=-1.7474e-13
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_14=-0.18283
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_14=-5.8145e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_14=0.043819
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_14=-0.0003715
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_14=-0.084668
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_14=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_14=-5.06e-11
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_15=-0.10493
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_15=-0.0066134
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_15=-0.36319
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_15=-3.1989e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_15=-0.19516
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_15=-1.1952e-18
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_15=-0.0011793
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_15=-12316.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_15=-4.5e-7
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_15=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_16=-7.4858e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_16=-0.046726
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_16=-0.0029649
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_16=0.10812
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_16=5.1967e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_16=-0.14571
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_16=-2.5784e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_16=0.037966
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_16=-0.0027377
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_16=-1.3973e-6
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_16=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_16=-0.10779
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_17=-0.0074577
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_17=-0.04734
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_17=1.8017e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_17=-0.036843
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_17=-0.012322
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_17=0.21238
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_17=3.4276e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_17=-0.24376
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_17=-2.2984e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_17=0.0074847
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_17=-0.0021369
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_17=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_18=-0.0019436
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_18=-0.08591
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_18=-0.015327
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_18=3.542e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_18=-0.025337
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_18=-0.016989
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_18=0.38189
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_18=2.6195e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_18=-0.32122
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_18=-2.1799e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_18=0.0014114
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_18=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_19=-0.001547
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_19=-0.099999
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_19=-0.0093411
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_19=3.4023e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_19=-0.026846
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_19=-0.01926
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_19=0.6214
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_19=2.6177e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_19=-0.38313
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_19=-1.1567e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_19=0.00015762
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_20=-0.0008493
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_20=-11352.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_20=-0.1126
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_20=0.0013192
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_20=-0.15791
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_20=-0.25975
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_20=6.6964e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_20=2.9253e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_21=-0.00014915
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_21=-11412.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_21=1.0947e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_21=-0.060457
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_21=-0.0042354
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_21=-0.18888
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_21=-0.23
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_21=4.9625e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_21=3.3096e-19
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_22=-0.2219
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_22=-2.3943e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_22=0.032162
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_22=-0.0018579
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_22=-0.093515
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_22=-9.7177e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_22=-0.047547
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_22=0.0079029
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_22=-0.057691
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_22=1.9974e-12
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_23=0.10024
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_23=4.9398e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_23=-0.30353
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_23=-3.2795e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_23=0.00028143
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_23=-0.0030795
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_23=-0.0079285
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_23=-0.014367
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_23=-3.6886e-12
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_23=-0.033013
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_23=-0.0030642
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_24=-0.0067096
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_24=0.35211
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_24=4.2158e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_24=-0.30203
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_24=-4.0315e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_24=0.001735
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_24=-0.0031364
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_24=-0.078814
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_24=-0.013816
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_24=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_24=-8.8875e-14
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_24=-0.026086
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_25=-0.0208
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_25=-0.0098344
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_25=0.56435
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_25=4.1901e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_25=-0.3615
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_25=-3.0855e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_25=0.00053738
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_25=-0.0028418
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_25=-0.099951
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_25=-0.0054488
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_25=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_25=-2.5927e-13
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_26=-0.11131
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_26=-0.0055458
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_26=-0.28683
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_26=4.2929e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_26=-0.17933
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_26=2.7713e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_26=-3.6655e-5
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_26=-10490.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_26=3.0e-7
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_26=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_27=5.3028e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_27=-0.05027
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_27=0.0035792
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_27=-0.28192
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_27=2.7136e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_27=-0.24717
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_27=2.5526e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_27=0.00031269
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_27=-9644.7
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_27=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_28=3.3821e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_28=-0.051336
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_28=0.010605
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_28=-0.12
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_28=3.1807e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_28=-0.29105
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_28=-1.0796e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_28=-0.0013987
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_28=-9154.7
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_28=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_29=-0.0030942
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_29=-6.9772e-7
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_29=-0.092123
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_29=-5.06e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_29=-0.046661
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_29=0.0068682
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_29=0.084807
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_29=4.5534e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_29=-0.075506
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_29=-4.414e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_29=0.027943
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_29=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_30=-0.0038175
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_30=-0.0045198
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_30=-0.023244
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_30=-3.0162e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_30=-0.033692
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_30=-0.0031254
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_30=-0.14808
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_30=0.20267
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_30=5.2436e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_30=-5.357e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_30=0.0020451
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_31=0.0022363
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_31=-0.0032561
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_31=-0.064893
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_31=-0.016796
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_31=-1.2695e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_31=-0.027851
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_31=-0.0080288
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_31=-0.25424
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_31=0.25558
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_31=4.1919e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_31=-4.5483e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_32=-0.00033374
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_32=-0.0031495
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_32=-0.0063838
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_32=-1.3284e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_32=-0.023384
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_32=-0.0092581
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_32=-0.33806
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_32=0.99453
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_32=4.4861e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_32=-3.862e-19
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_33=-0.1868
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_33=3.1635e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_33=0.00076765
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_33=-8082.5
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_33=-0.11328
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_33=-0.0049124
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_33=-0.31419
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_33=2.5342e-12
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_34=-0.170321
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_34=3.4845e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_34=-0.27802
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_34=-4.3629e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_34=-0.0028047
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_34=-11258.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_34=1.0432e-11
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_34=-0.047284
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_34=0.0096808
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_35=-0.013148
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_35=0.1047
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_35=1.2125e-11
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_35=-0.083988
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_35=4.7539e-20
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_35=-0.003457
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_35=2.6925e-7
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_35=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_35=-2.4215e-9
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_35=2.1644e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_35=-0.12204
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_36=-0.058569
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_36=-0.01786
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_36=0.99372
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_36=6.4917e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_36=-0.53925
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_36=-1.8362e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_36=-0.003775
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_36=-0.1
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_36=5.9604e-8
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_36=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_36=4.2551e-10
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_36=4.3256e-10
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_37=3.3626e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_37=-0.066111
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_37=-0.019646
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_37=0.32331
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_37=7.1708e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_37=-0.23808
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_37=-1.1404e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_37=-0.0026716
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_37=9.5177e-8
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_37=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_37=-1.5823e-9
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_38=-3.398e-9
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_38=4.4079e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_38=-0.068451
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_38=-0.016156
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_38=0.34571
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_38=1.0732e-11
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_38=-0.42153
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_38=-1.6411e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_38=-0.0042034
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_38=4.885e-8
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_38=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_39=5.7403e-8
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_39=3.3719e-8
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_39=4.4337e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_39=-0.064273
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_39=-0.02017
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_39=0.52754
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_39=8.1318e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_39=-0.56147
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_39=-3.653e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_39=-0.0041811
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_39=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_40=8.06e-10
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_40=-0.15277
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_40=0.0011713
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_40=-0.18048
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_40=-0.13975
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_40=3.7351e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_40=2.2029e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_40=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_40=-0.0027234
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_40=-23997.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_41=-0.0025844
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_41=-21982.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_41=6.9406e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_41=-0.13143
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_41=-0.015942
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_41=-0.07378
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_41=-0.13088863
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_41=3.912e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_41=3.6155e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_41=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_42=-0.0021575
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_42=-17815.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_42=8.06e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_42=-0.1381
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_42=-0.022906
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_42=-0.1599
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_42=1.2974e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_42=1.7324e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_42=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_43=-0.0015022
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_43=2.5083e-7
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_43=1.8595e-9
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_43=1.5619e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_43=-0.057516
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_43=-0.00361
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_43=-0.11492
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_43=0.15731
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_43=5.6688e-12
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_43=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_43=9.2328e-20
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_44=-0.23784
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_44=1.4394e-20
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_44=-0.001027
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_44=1.2039e-7
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_44=-2.0663e-10
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_44=2.0984e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_44=-0.062774
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_44=-0.013153
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_44=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_44=0.32388
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_44=3.7152e-12
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_45=0.34189
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_45=2.6165e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_45=-0.42112
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_45=-2.3003e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_45=-0.0020521
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_45=1.597e-7
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_45=-1.606e-10
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_45=2.5642e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_45=-0.038017
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_45=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_45=-0.018074
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_46=0.0035731
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_46=-0.100982
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_46=1.293e-11
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_46=-0.17395
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_46=6.3502e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_46=-0.001157
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_46=-17789.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_46=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_46=8.06e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_46=-0.13699
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_47=-0.065441
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_47=-0.00085911
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_47=0.12718
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_47=4.9518e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_47=-0.12752
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_47=8.6671e-20
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_47=-0.0011573
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_47=-17521.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_47=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_47=2.9655e-10
.param sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_48=4.6959e-10
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_48=-0.099532
.param sky130_fd_pr__nfet_g5v0d10v5__keta_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__k2_diff_48=5.4148e-5
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_48=-0.05129
.param sky130_fd_pr__nfet_g5v0d10v5__ua_diff_48=8.8919e-12
.param sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_48=-0.092595
.param sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ub_diff_48=2.3132e-19
.param sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__a0_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__u0_diff_48=-0.0018033
.param sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_48=-20000.0
.param sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b0_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__ags_diff_48=0.0
.param sky130_fd_pr__nfet_g5v0d10v5__b1_diff_48=0.0
.include "sky130_fd_pr__nfet_g5v0d10v5.pm3.spice"