* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_03v3_nvt__toxe_mult=0.9635
.param sky130_fd_pr__nfet_03v3_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_03v3_nvt__overlap_mult=0.51025
.param sky130_fd_pr__nfet_03v3_nvt__ajunction_mult=0.68772
.param sky130_fd_pr__nfet_03v3_nvt__pjunction_mult=0.9019
.param sky130_fd_pr__nfet_03v3_nvt__lint_diff=1.21275e-8
.param sky130_fd_pr__nfet_03v3_nvt__wint_diff=-2.252e-8
.param sky130_fd_pr__nfet_03v3_nvt__dlc_diff=1.6112e-8
.param sky130_fd_pr__nfet_03v3_nvt__dwc_diff=-2.252e-8
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_0=0.017139
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_0=-0.016856
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_0=-1.0949
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_0=-0.041263
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_0=0.00079908
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_0=-1877.8
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_0=-8.8355e-20
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_0=1.2237e-11
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_1=3.5287e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_1=0.010252
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_1=-0.00051272
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_1=-1.3847
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_1=-0.0485
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_1=-7.0468e-5
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_1=-9793.6
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_1=2.2579e-19
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_2=1.2013e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_2=1.1421e-10
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_2=0.0012159
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_2=-0.49031
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_2=-0.034235
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_2=0.0043842
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_2=-8139.1
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_3=6.5751e-20
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_3=2.2944e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_3=0.0177
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_3=-0.01428
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_3=-1.0283
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_3=-0.04376
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_3=0.0014903
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_3=-3761.4
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_4=-4.2142e-19
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_4=-1.3052e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_4=0.044934
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_4=0.0083971
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_4=-1.5502
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_4=-0.068861
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_4=0.0016304
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_4=-6110.3
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_5=0.01509
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_5=-5015.2
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_5=2.0257e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_5=4.4064e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_5=0.0059498
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_5=-1.6314
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_5=0.014604
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_6=-0.77252
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_6=-0.0039098
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_6=0.011371
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_6=-3438.4
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_6=1.7785e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_6=5.037e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_6=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_6=0.0058775
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_7=0.021791
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_7=0.0022917
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_7=-1.3041
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_7=-0.046002
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_7=0.00087134
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_7=-9538.4
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_7=4.1235e-19
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_7=2.4503e-11
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_03v3_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__b0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__k2_diff_8=0.0038297
.param sky130_fd_pr__nfet_03v3_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__nfactor_diff_8=-0.51817
.param sky130_fd_pr__nfet_03v3_nvt__vth0_diff_8=-0.040702
.param sky130_fd_pr__nfet_03v3_nvt__u0_diff_8=0.006163
.param sky130_fd_pr__nfet_03v3_nvt__vsat_diff_8=-7789.7
.param sky130_fd_pr__nfet_03v3_nvt__b1_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ub_diff_8=1.381e-18
.param sky130_fd_pr__nfet_03v3_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__ua_diff_8=1.3573e-10
.param sky130_fd_pr__nfet_03v3_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_03v3_nvt__pclm_diff_8=0.0
.include "sky130_fd_pr__nfet_03v3_nvt.pm3.spice"