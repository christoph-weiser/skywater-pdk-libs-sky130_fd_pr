* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8__toxe_mult=0.9635
.param sky130_fd_pr__nfet_01v8__rshn_mult=1.0
.param sky130_fd_pr__nfet_01v8__overlap_mult=0.95013
.param sky130_fd_pr__nfet_01v8__lint_diff=1.21275e-8
.param sky130_fd_pr__nfet_01v8__wint_diff=-2.252e-8
.param sky130_fd_pr__nfet_01v8__dlc_diff=8.0874e-9
.param sky130_fd_pr__nfet_01v8__dwc_diff=-2.252e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_0=-1.8425e-19
.param sky130_fd_pr__nfet_01v8__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_0=5.685e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_0=-29297.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_0=0.041243
.param sky130_fd_pr__nfet_01v8__vth0_diff_0=-0.10074
.param sky130_fd_pr__nfet_01v8__nfactor_diff_0=0.8236
.param sky130_fd_pr__nfet_01v8__u0_diff_0=-0.005854
.param sky130_fd_pr__nfet_01v8__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_0=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_1=-1.3801e-19
.param sky130_fd_pr__nfet_01v8__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_1=4.7162e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_1=-22217.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_1=0.039934
.param sky130_fd_pr__nfet_01v8__vth0_diff_1=-0.069738
.param sky130_fd_pr__nfet_01v8__nfactor_diff_1=0.85772
.param sky130_fd_pr__nfet_01v8__u0_diff_1=-0.0049428
.param sky130_fd_pr__nfet_01v8__nfactor_diff_2=1.1356
.param sky130_fd_pr__nfet_01v8__u0_diff_2=0.0013905
.param sky130_fd_pr__nfet_01v8__vth0_diff_2=-0.0020947
.param sky130_fd_pr__nfet_01v8__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_2=2.6748e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_2=-2.9823e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_2=-0.07434
.param sky130_fd_pr__nfet_01v8__a0_diff_2=0.30304
.param sky130_fd_pr__nfet_01v8__b0_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_2=-0.0053077
.param sky130_fd_pr__nfet_01v8__keta_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_3=-0.0046106
.param sky130_fd_pr__nfet_01v8__nfactor_diff_3=0.84258
.param sky130_fd_pr__nfet_01v8__u0_diff_3=0.00078603
.param sky130_fd_pr__nfet_01v8__vth0_diff_3=-0.0087266
.param sky130_fd_pr__nfet_01v8__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_3=2.3573e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_3=-1.6853e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_3=-0.032489
.param sky130_fd_pr__nfet_01v8__a0_diff_3=0.067824
.param sky130_fd_pr__nfet_01v8__b0_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_4=0.0041217
.param sky130_fd_pr__nfet_01v8__nfactor_diff_4=1.0497
.param sky130_fd_pr__nfet_01v8__u0_diff_4=-0.00092253
.param sky130_fd_pr__nfet_01v8__vth0_diff_4=-0.012158
.param sky130_fd_pr__nfet_01v8__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_4=1.0247e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_4=3.5347e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_4=-0.0078262
.param sky130_fd_pr__nfet_01v8__a0_diff_4=0.023077
.param sky130_fd_pr__nfet_01v8__b0_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_5=0.0058164
.param sky130_fd_pr__nfet_01v8__nfactor_diff_5=0.88776
.param sky130_fd_pr__nfet_01v8__u0_diff_5=-0.0010888
.param sky130_fd_pr__nfet_01v8__vth0_diff_5=-0.0096783
.param sky130_fd_pr__nfet_01v8__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_5=1.0006e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_5=4.0462e-12
.param sky130_fd_pr__nfet_01v8__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_5=-0.016825
.param sky130_fd_pr__nfet_01v8__a0_diff_5=0.034496
.param sky130_fd_pr__nfet_01v8__b0_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_6=0.039149
.param sky130_fd_pr__nfet_01v8__nfactor_diff_6=1.309
.param sky130_fd_pr__nfet_01v8__u0_diff_6=-0.0059282
.param sky130_fd_pr__nfet_01v8__vth0_diff_6=-0.082368
.param sky130_fd_pr__nfet_01v8__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_6=-2.5891e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_6=5.5593e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_6=-30394.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_6=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_7=0.022032
.param sky130_fd_pr__nfet_01v8__nfactor_diff_7=0.63926
.param sky130_fd_pr__nfet_01v8__u0_diff_7=-0.0033503
.param sky130_fd_pr__nfet_01v8__vth0_diff_7=-0.061613
.param sky130_fd_pr__nfet_01v8__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_7=-2.4572e-20
.param sky130_fd_pr__nfet_01v8__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_7=3.4046e-11
.param sky130_fd_pr__nfet_01v8__vsat_diff_7=-28245.0
.param sky130_fd_pr__nfet_01v8__a0_diff_7=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_8=1.9021e-11
.param sky130_fd_pr__nfet_01v8__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_8=0.0076402
.param sky130_fd_pr__nfet_01v8__nfactor_diff_8=1.3774
.param sky130_fd_pr__nfet_01v8__u0_diff_8=-0.0012732
.param sky130_fd_pr__nfet_01v8__vth0_diff_8=-0.037767
.param sky130_fd_pr__nfet_01v8__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_8=2.9793e-19
.param sky130_fd_pr__nfet_01v8__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_8=-28984.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_9=-2.7776e-20
.param sky130_fd_pr__nfet_01v8__vsat_diff_9=-17190.0
.param sky130_fd_pr__nfet_01v8__a0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_9=7.254e-12
.param sky130_fd_pr__nfet_01v8__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_9=0.0057044
.param sky130_fd_pr__nfet_01v8__nfactor_diff_9=1.4725
.param sky130_fd_pr__nfet_01v8__u0_diff_9=-0.0021368
.param sky130_fd_pr__nfet_01v8__vth0_diff_9=-0.0074743
.param sky130_fd_pr__nfet_01v8__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_9=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_10=0.04236
.param sky130_fd_pr__nfet_01v8__ua_diff_10=4.1917e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_10=-1.4028e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_10=-26960.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_10=-0.064685
.param sky130_fd_pr__nfet_01v8__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_10=0.94373
.param sky130_fd_pr__nfet_01v8__u0_diff_10=-0.0043223
.param sky130_fd_pr__nfet_01v8__pclm_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_11=0.90212
.param sky130_fd_pr__nfet_01v8__u0_diff_11=0.00025182
.param sky130_fd_pr__nfet_01v8__ags_diff_11=-0.04068
.param sky130_fd_pr__nfet_01v8__keta_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_11=-0.0018907
.param sky130_fd_pr__nfet_01v8__ua_diff_11=-6.8936e-13
.param sky130_fd_pr__nfet_01v8__eta0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_11=1.3995e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_11=0.013802
.param sky130_fd_pr__nfet_01v8__rdsw_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_11=0.0030064
.param sky130_fd_pr__nfet_01v8__pdits_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_11=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_12=1.0365
.param sky130_fd_pr__nfet_01v8__u0_diff_12=-0.0023921
.param sky130_fd_pr__nfet_01v8__ags_diff_12=0.0048249
.param sky130_fd_pr__nfet_01v8__keta_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_12=0.002976
.param sky130_fd_pr__nfet_01v8__ua_diff_12=7.4962e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_12=-8.8622e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_12=0.013456
.param sky130_fd_pr__nfet_01v8__rdsw_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_12=-0.010504
.param sky130_fd_pr__nfet_01v8__pdits_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_12=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_13=1.3067
.param sky130_fd_pr__nfet_01v8__u0_diff_13=-0.0033083
.param sky130_fd_pr__nfet_01v8__ags_diff_13=0.030222
.param sky130_fd_pr__nfet_01v8__keta_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_13=0.0045206
.param sky130_fd_pr__nfet_01v8__ua_diff_13=1.8203e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_13=-1.8415e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_13=-0.018323
.param sky130_fd_pr__nfet_01v8__rdsw_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_13=-0.011631
.param sky130_fd_pr__nfet_01v8__b0_diff_13=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_14=1.0962
.param sky130_fd_pr__nfet_01v8__u0_diff_14=-0.0023253
.param sky130_fd_pr__nfet_01v8__ags_diff_14=0.0051407
.param sky130_fd_pr__nfet_01v8__keta_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_14=0.0058036
.param sky130_fd_pr__nfet_01v8__ua_diff_14=6.5432e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_14=-1.2092e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_14=0.016324
.param sky130_fd_pr__nfet_01v8__rdsw_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_14=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_14=-0.0078698
.param sky130_fd_pr__nfet_01v8__kt1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_15=-22922.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_15=-0.08669
.param sky130_fd_pr__nfet_01v8__b0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_15=1.1095
.param sky130_fd_pr__nfet_01v8__u0_diff_15=-0.0070567
.param sky130_fd_pr__nfet_01v8__ags_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_15=0.048668
.param sky130_fd_pr__nfet_01v8__ua_diff_15=5.684e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_15=-5.3557e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_15=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_16=-20211.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_16=-0.043878
.param sky130_fd_pr__nfet_01v8__b0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_16=0.5721
.param sky130_fd_pr__nfet_01v8__u0_diff_16=-0.0030356
.param sky130_fd_pr__nfet_01v8__ags_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_16=0.033098
.param sky130_fd_pr__nfet_01v8__ua_diff_16=3.0616e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_16=-2.118e-21
.param sky130_fd_pr__nfet_01v8__tvoff_diff_16=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_17=-19092.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_17=-0.034533
.param sky130_fd_pr__nfet_01v8__pdits_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_17=1.2421
.param sky130_fd_pr__nfet_01v8__u0_diff_17=-0.00041085
.param sky130_fd_pr__nfet_01v8__ags_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_17=0.015329
.param sky130_fd_pr__nfet_01v8__ua_diff_17=6.6214e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_17=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_17=1.6031e-19
.param sky130_fd_pr__nfet_01v8__ub_diff_18=1.032e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_18=-4614.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_18=-0.014924
.param sky130_fd_pr__nfet_01v8__pdits_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_18=0.9249
.param sky130_fd_pr__nfet_01v8__u0_diff_18=-0.0011111
.param sky130_fd_pr__nfet_01v8__ags_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_18=0.0043522
.param sky130_fd_pr__nfet_01v8__ua_diff_18=4.3593e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_18=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__ua_diff_19=-3.7829e-14
.param sky130_fd_pr__nfet_01v8__ub_diff_19=1.2662e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_19=0.026691
.param sky130_fd_pr__nfet_01v8__rdsw_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_19=0.0027493
.param sky130_fd_pr__nfet_01v8__pdits_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_19=0.85527
.param sky130_fd_pr__nfet_01v8__u0_diff_19=-9.7139e-5
.param sky130_fd_pr__nfet_01v8__ags_diff_19=0.061189
.param sky130_fd_pr__nfet_01v8__keta_diff_19=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_19=0.004984
.param sky130_fd_pr__nfet_01v8__ua_diff_20=1.1526e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_20=-2.4487e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_20=-0.0027531
.param sky130_fd_pr__nfet_01v8__rdsw_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_20=-0.014574
.param sky130_fd_pr__nfet_01v8__pdits_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_20=0.99163
.param sky130_fd_pr__nfet_01v8__u0_diff_20=-0.0036938
.param sky130_fd_pr__nfet_01v8__ags_diff_20=0.018914
.param sky130_fd_pr__nfet_01v8__keta_diff_20=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_20=0.0030348
.param sky130_fd_pr__nfet_01v8__ags_diff_21=-0.015591
.param sky130_fd_pr__nfet_01v8__keta_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_21=0.0025752
.param sky130_fd_pr__nfet_01v8__ua_diff_21=6.8301e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_21=-1.5459e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_21=0.032179
.param sky130_fd_pr__nfet_01v8__rdsw_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_21=-0.010241
.param sky130_fd_pr__nfet_01v8__pdits_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_21=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_21=0.82101
.param sky130_fd_pr__nfet_01v8__u0_diff_21=-0.0022896
.param sky130_fd_pr__nfet_01v8__pclm_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_22=1.0794
.param sky130_fd_pr__nfet_01v8__u0_diff_22=-0.0015731
.param sky130_fd_pr__nfet_01v8__ags_diff_22=0.031797
.param sky130_fd_pr__nfet_01v8__keta_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_22=0.0062222
.param sky130_fd_pr__nfet_01v8__ua_diff_22=4.5017e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_22=-4.929e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_22=-0.018961
.param sky130_fd_pr__nfet_01v8__rdsw_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_22=-0.0052112
.param sky130_fd_pr__nfet_01v8__pdits_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_22=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_23=1.4808
.param sky130_fd_pr__nfet_01v8__u0_diff_23=-0.0023173
.param sky130_fd_pr__nfet_01v8__ags_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_23=0.040162
.param sky130_fd_pr__nfet_01v8__ua_diff_23=1.6728e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_23=-7.9157e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_23=-16743.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_23=-0.069697
.param sky130_fd_pr__nfet_01v8__pdits_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_23=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_24=1.5509
.param sky130_fd_pr__nfet_01v8__u0_diff_24=-0.0095729
.param sky130_fd_pr__nfet_01v8__ags_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_24=0.03105
.param sky130_fd_pr__nfet_01v8__ua_diff_24=7.8244e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_24=-5.4162e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_24=-15248.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_24=-0.061307
.param sky130_fd_pr__nfet_01v8__b0_diff_24=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_25=1.0158
.param sky130_fd_pr__nfet_01v8__u0_diff_25=-0.00030254
.param sky130_fd_pr__nfet_01v8__ags_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_25=0.013824
.param sky130_fd_pr__nfet_01v8__ua_diff_25=6.2221e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_25=1.8421e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_25=-16202.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_25=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_25=-0.017264
.param sky130_fd_pr__nfet_01v8__kt1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_26=-7360.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_26=-0.010605
.param sky130_fd_pr__nfet_01v8__b0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_26=1.0973
.param sky130_fd_pr__nfet_01v8__u0_diff_26=-0.00075949
.param sky130_fd_pr__nfet_01v8__ags_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_26=0.002474
.param sky130_fd_pr__nfet_01v8__ua_diff_26=2.3906e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_26=3.4242e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_26=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_27=0.025136
.param sky130_fd_pr__nfet_01v8__rdsw_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_27=-0.012606
.param sky130_fd_pr__nfet_01v8__b0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_27=0.94796
.param sky130_fd_pr__nfet_01v8__u0_diff_27=-0.0012564
.param sky130_fd_pr__nfet_01v8__ags_diff_27=-0.01694
.param sky130_fd_pr__nfet_01v8__keta_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_27=0.0034005
.param sky130_fd_pr__nfet_01v8__ua_diff_27=4.7202e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_27=3.6896e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_27=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_28=-0.025217
.param sky130_fd_pr__nfet_01v8__rdsw_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_28=-0.0054922
.param sky130_fd_pr__nfet_01v8__pdits_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_28=0.92951
.param sky130_fd_pr__nfet_01v8__u0_diff_28=-0.0011803
.param sky130_fd_pr__nfet_01v8__ags_diff_28=0.03232
.param sky130_fd_pr__nfet_01v8__keta_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_28=0.0042396
.param sky130_fd_pr__nfet_01v8__ua_diff_28=4.0266e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_28=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_28=1.4013e-20
.param sky130_fd_pr__nfet_01v8__ub_diff_29=5.3622e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_29=-0.057732
.param sky130_fd_pr__nfet_01v8__rdsw_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_29=-0.0085008
.param sky130_fd_pr__nfet_01v8__pdits_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_29=0.83848
.param sky130_fd_pr__nfet_01v8__u0_diff_29=-0.00077347
.param sky130_fd_pr__nfet_01v8__ags_diff_29=0.047346
.param sky130_fd_pr__nfet_01v8__keta_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_29=0.002189
.param sky130_fd_pr__nfet_01v8__ua_diff_29=2.8611e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_29=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_30=-1.8733e-21
.param sky130_fd_pr__nfet_01v8__tvoff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_30=-0.023064
.param sky130_fd_pr__nfet_01v8__rdsw_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_30=-0.00010044
.param sky130_fd_pr__nfet_01v8__pdits_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_30=0.78189
.param sky130_fd_pr__nfet_01v8__u0_diff_30=-0.00069527
.param sky130_fd_pr__nfet_01v8__ags_diff_30=0.031119
.param sky130_fd_pr__nfet_01v8__keta_diff_30=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_30=0.0042181
.param sky130_fd_pr__nfet_01v8__ua_diff_30=1.9583e-12
.param sky130_fd_pr__nfet_01v8__ua_diff_31=4.1896e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_31=2.0152e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_31=-12204.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_31=-0.048836
.param sky130_fd_pr__nfet_01v8__pdits_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_31=-0.11472
.param sky130_fd_pr__nfet_01v8__u0_diff_31=0.00050692
.param sky130_fd_pr__nfet_01v8__ags_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_31=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_31=0.034176
.param sky130_fd_pr__nfet_01v8__ags_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_32=0.029531
.param sky130_fd_pr__nfet_01v8__ua_diff_32=6.8335e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_32=-4.0465e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_32=-14690.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_32=-0.053486
.param sky130_fd_pr__nfet_01v8__pdits_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_32=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_32=1.4435
.param sky130_fd_pr__nfet_01v8__u0_diff_32=-0.0079835
.param sky130_fd_pr__nfet_01v8__pclm_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_33=0.75301
.param sky130_fd_pr__nfet_01v8__u0_diff_33=-0.00044388
.param sky130_fd_pr__nfet_01v8__ags_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_33=0.014786
.param sky130_fd_pr__nfet_01v8__ua_diff_33=6.4858e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_33=1.3291e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_33=-17397.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_33=-0.017301
.param sky130_fd_pr__nfet_01v8__pdits_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_33=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_34=1.0269
.param sky130_fd_pr__nfet_01v8__u0_diff_34=-0.0007785
.param sky130_fd_pr__nfet_01v8__ags_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_34=0.0023824
.param sky130_fd_pr__nfet_01v8__ua_diff_34=2.4627e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_34=3.1021e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_34=-5303.6
.param sky130_fd_pr__nfet_01v8__kt1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_34=-0.012707
.param sky130_fd_pr__nfet_01v8__pdits_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_34=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_35=9.3829e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_35=2.1945
.param sky130_fd_pr__nfet_01v8__u0_diff_35=-0.002626
.param sky130_fd_pr__nfet_01v8__ags_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_35=0.0024195
.param sky130_fd_pr__nfet_01v8__ua_diff_35=8.799e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_35=7.7707e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_35=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_35=-0.034885
.param sky130_fd_pr__nfet_01v8__b0_diff_35=-3.549e-8
.param sky130_fd_pr__nfet_01v8__b0_diff_36=6.3469e-8
.param sky130_fd_pr__nfet_01v8__pdits_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_36=2.5194e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_36=1.0826
.param sky130_fd_pr__nfet_01v8__u0_diff_36=-0.0013127
.param sky130_fd_pr__nfet_01v8__ags_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_36=0.0018953
.param sky130_fd_pr__nfet_01v8__ua_diff_36=3.9032e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_36=8.9052e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_36=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_36=-0.0048969
.param sky130_fd_pr__nfet_01v8__kt1_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_37=-0.056501
.param sky130_fd_pr__nfet_01v8__b0_diff_37=1.3378e-7
.param sky130_fd_pr__nfet_01v8__pdits_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_37=6.8667e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_37=1.6485
.param sky130_fd_pr__nfet_01v8__u0_diff_37=-0.003765
.param sky130_fd_pr__nfet_01v8__ags_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_37=0.0042254
.param sky130_fd_pr__nfet_01v8__ua_diff_37=1.2314e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_37=-4.279e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_37=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_38=-0.035395
.param sky130_fd_pr__nfet_01v8__b0_diff_38=6.1085e-8
.param sky130_fd_pr__nfet_01v8__pdits_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_38=8.4199e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_38=1.2757
.param sky130_fd_pr__nfet_01v8__u0_diff_38=-0.0022926
.param sky130_fd_pr__nfet_01v8__ags_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_38=0.0090756
.param sky130_fd_pr__nfet_01v8__ua_diff_38=7.918e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_38=9.0819e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_38=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_39=-0.0056917
.param sky130_fd_pr__nfet_01v8__pdits_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_39=7.9741e-8
.param sky130_fd_pr__nfet_01v8__b1_diff_39=2.1557e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_39=0.9785
.param sky130_fd_pr__nfet_01v8__u0_diff_39=-0.0016882
.param sky130_fd_pr__nfet_01v8__ags_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_39=-0.0015846
.param sky130_fd_pr__nfet_01v8__ua_diff_39=5.052e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_39=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_39=4.2656e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_40=-42474.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_40=-0.14746
.param sky130_fd_pr__nfet_01v8__pdits_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_40=1.0604
.param sky130_fd_pr__nfet_01v8__u0_diff_40=-0.0066881
.param sky130_fd_pr__nfet_01v8__ags_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_40=0.034077
.param sky130_fd_pr__nfet_01v8__ua_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_40=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_41=1.0874e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_41=-45699.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_41=-0.10449
.param sky130_fd_pr__nfet_01v8__pdits_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_41=0.98392
.param sky130_fd_pr__nfet_01v8__u0_diff_41=-0.0055054
.param sky130_fd_pr__nfet_01v8__ags_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_41=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_41=0.0088642
.param sky130_fd_pr__nfet_01v8__ua_diff_41=3.1502e-11
.param sky130_fd_pr__nfet_01v8__ua_diff_42=1.0002e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_42=1.0334e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_42=-51798.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_42=-0.029837
.param sky130_fd_pr__nfet_01v8__pdits_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_42=1.6886
.param sky130_fd_pr__nfet_01v8__u0_diff_42=-0.0025307
.param sky130_fd_pr__nfet_01v8__ags_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_42=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_42=0.0082221
.param sky130_fd_pr__nfet_01v8__ags_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_43=0.0094379
.param sky130_fd_pr__nfet_01v8__ua_diff_43=1.2467e-13
.param sky130_fd_pr__nfet_01v8__eta0_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_43=2.5516e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_43=-0.014814
.param sky130_fd_pr__nfet_01v8__pdits_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_43=1.9371e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_43=6.2753e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_43=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_43=1.8005
.param sky130_fd_pr__nfet_01v8__u0_diff_43=0.00012802
.param sky130_fd_pr__nfet_01v8__pclm_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_44=1.4439
.param sky130_fd_pr__nfet_01v8__u0_diff_44=-0.0054279
.param sky130_fd_pr__nfet_01v8__ags_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_44=0.0041381
.param sky130_fd_pr__nfet_01v8__ua_diff_44=1.603e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_44=-2.6649e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_44=-0.032691
.param sky130_fd_pr__nfet_01v8__pdits_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_44=1.3999e-7
.param sky130_fd_pr__nfet_01v8__voff_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_44=8.5735e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_44=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_45=1.3136
.param sky130_fd_pr__nfet_01v8__u0_diff_45=-0.002825
.param sky130_fd_pr__nfet_01v8__ags_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_45=0.0044471
.param sky130_fd_pr__nfet_01v8__ua_diff_45=8.6251e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_45=-3.8973e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_45=-0.017554
.param sky130_fd_pr__nfet_01v8__pdits_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_45=9.4644e-8
.param sky130_fd_pr__nfet_01v8__voff_diff_45=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_45=4.0028e-9
.param sky130_fd_pr__nfet_01v8__pdits_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_46=1.5919e-9
.param sky130_fd_pr__nfet_01v8__pditsd_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_46=0.71682
.param sky130_fd_pr__nfet_01v8__u0_diff_46=-0.00086513
.param sky130_fd_pr__nfet_01v8__ags_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_46=0.0023491
.param sky130_fd_pr__nfet_01v8__ua_diff_46=3.625e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_46=1.6356e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_46=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_46=-0.0040694
.param sky130_fd_pr__nfet_01v8__b0_diff_46=6.024e-8
.param sky130_fd_pr__nfet_01v8__b0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_47=0.99292
.param sky130_fd_pr__nfet_01v8__u0_diff_47=-0.0065314
.param sky130_fd_pr__nfet_01v8__ags_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_47=0.033937
.param sky130_fd_pr__nfet_01v8__ua_diff_47=3.5207e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_47=-2.7169e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_47=-44229.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_47=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_47=-0.13487
.param sky130_fd_pr__nfet_01v8__kt1_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_48=-40596.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_48=-0.031371
.param sky130_fd_pr__nfet_01v8__b0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_48=1.6077
.param sky130_fd_pr__nfet_01v8__u0_diff_48=-0.00011217
.param sky130_fd_pr__nfet_01v8__ags_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_48=0.0020322
.param sky130_fd_pr__nfet_01v8__ua_diff_48=7.8961e-12
.param sky130_fd_pr__nfet_01v8__eta0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_48=1.9998e-19
.param sky130_fd_pr__nfet_01v8__tvoff_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_48=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_49=-29107.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_49=-0.083391
.param sky130_fd_pr__nfet_01v8__b0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_49=0.80364
.param sky130_fd_pr__nfet_01v8__u0_diff_49=-0.0038179
.param sky130_fd_pr__nfet_01v8__ags_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_49=0.03982
.param sky130_fd_pr__nfet_01v8__ua_diff_49=4.0178e-11
.param sky130_fd_pr__nfet_01v8__eta0_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_49=6.7996e-20
.param sky130_fd_pr__nfet_01v8__tvoff_diff_49=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_50=-29827.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_50=-0.10606
.param sky130_fd_pr__nfet_01v8__pdits_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__nfactor_diff_50=0.56382
.param sky130_fd_pr__nfet_01v8__u0_diff_50=-0.0050668
.param sky130_fd_pr__nfet_01v8__ags_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__keta_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_50=0.035186
.param sky130_fd_pr__nfet_01v8__ua_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__eta0_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__ub_diff_50=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_51=-33982.49122578
.param sky130_fd_pr__nfet_01v8__kt1_diff_51=4.36291e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_51=-0.0912518
.param sky130_fd_pr__nfet_01v8__pdits_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_51=0.00023948
.param sky130_fd_pr__nfet_01v8__u0_diff_51=-0.00172097
.param sky130_fd_pr__nfet_01v8__nfactor_diff_51=0.28498727
.param sky130_fd_pr__nfet_01v8__keta_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_51=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_51=0.03496439
.param sky130_fd_pr__nfet_01v8__ua_diff_51=6.38272e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_51=8.82259e-20
.param sky130_fd_pr__nfet_01v8__eta0_diff_51=-2.08167e-17
.param sky130_fd_pr__nfet_01v8__ub_diff_52=-9.88831e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_52=2.39904e-5
.param sky130_fd_pr__nfet_01v8__tvoff_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_52=-41493.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_52=-0.12103
.param sky130_fd_pr__nfet_01v8__pdits_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_52=0.0006774
.param sky130_fd_pr__nfet_01v8__u0_diff_52=-0.017441
.param sky130_fd_pr__nfet_01v8__nfactor_diff_52=0.32359691
.param sky130_fd_pr__nfet_01v8__keta_diff_52=0.00226031
.param sky130_fd_pr__nfet_01v8__ags_diff_52=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_52=0.029744
.param sky130_fd_pr__nfet_01v8__ua_diff_52=-1.6427e-12
.param sky130_fd_pr__nfet_01v8__ua_diff_53=2.59392e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_53=-8.07338e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_53=8.51883e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_53=-39855.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_53=-0.12287
.param sky130_fd_pr__nfet_01v8__pdits_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_53=0.00024054
.param sky130_fd_pr__nfet_01v8__u0_diff_53=-0.014549
.param sky130_fd_pr__nfet_01v8__nfactor_diff_53=0.32663125
.param sky130_fd_pr__nfet_01v8__keta_diff_53=0.00080262
.param sky130_fd_pr__nfet_01v8__ags_diff_53=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_53=0.029369
.param sky130_fd_pr__nfet_01v8__keta_diff_54=-0.00027377
.param sky130_fd_pr__nfet_01v8__ags_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_54=0.030064
.param sky130_fd_pr__nfet_01v8__ua_diff_54=1.64639e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_54=-2.86662e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_54=-2.90569e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_54=-41870.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_54=-0.13092
.param sky130_fd_pr__nfet_01v8__pdits_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_54=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_54=-8.20469e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_54=-0.0022189
.param sky130_fd_pr__nfet_01v8__nfactor_diff_54=0.35136061
.param sky130_fd_pr__nfet_01v8__pclm_diff_55=-3.03325e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_55=-0.0019602
.param sky130_fd_pr__nfet_01v8__nfactor_diff_55=0.35549327
.param sky130_fd_pr__nfet_01v8__keta_diff_55=-0.00010121
.param sky130_fd_pr__nfet_01v8__ags_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_55=0.030831
.param sky130_fd_pr__nfet_01v8__ua_diff_55=1.81079e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_55=-2.30916e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_55=-1.07421e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_55=-41866.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_55=-0.12602
.param sky130_fd_pr__nfet_01v8__pdits_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_55=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_56=-5.66337e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_56=0.00031229
.param sky130_fd_pr__nfet_01v8__nfactor_diff_56=0.34932529
.param sky130_fd_pr__nfet_01v8__keta_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_56=0.031119
.param sky130_fd_pr__nfet_01v8__ua_diff_56=2.25094e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_56=-5.55536e-20
.param sky130_fd_pr__nfet_01v8__eta0_diff_56=2.00573e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_56=-40931.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_56=-2.88948e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_56=-0.12242
.param sky130_fd_pr__nfet_01v8__pdits_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_56=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_57=-5.86462e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_57=0.0014122
.param sky130_fd_pr__nfet_01v8__nfactor_diff_57=0.34402866
.param sky130_fd_pr__nfet_01v8__keta_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_57=0.031396
.param sky130_fd_pr__nfet_01v8__ua_diff_57=2.47125e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_57=3.51976e-20
.param sky130_fd_pr__nfet_01v8__eta0_diff_57=2.077e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_57=-41388.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_57=-2.99216e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_57=-0.11936
.param sky130_fd_pr__nfet_01v8__b0_diff_57=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_58=-5.10014e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_58=0.0016098
.param sky130_fd_pr__nfet_01v8__nfactor_diff_58=0.34143761
.param sky130_fd_pr__nfet_01v8__keta_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_58=0.031526
.param sky130_fd_pr__nfet_01v8__ua_diff_58=2.57578e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_58=7.82369e-20
.param sky130_fd_pr__nfet_01v8__eta0_diff_58=1.80626e-6
.param sky130_fd_pr__nfet_01v8__tvoff_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_58=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_58=-41364.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_58=-2.60212e-5
.param sky130_fd_pr__nfet_01v8__vth0_diff_58=-0.11848
.param sky130_fd_pr__nfet_01v8__kt1_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_59=-33732.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_59=-0.1169
.param sky130_fd_pr__nfet_01v8__b0_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pdits_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_59=5.94765e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_59=0.0020456
.param sky130_fd_pr__nfet_01v8__nfactor_diff_59=0.32842233
.param sky130_fd_pr__nfet_01v8__keta_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_59=0.031651
.param sky130_fd_pr__nfet_01v8__ua_diff_59=2.61524e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_59=1.86252e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_59=-3.33296e-17
.param sky130_fd_pr__nfet_01v8__tvoff_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_59=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_60=-31573.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_60=-0.078715
.param sky130_fd_pr__nfet_01v8__pdits_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_60=5.9476e-5
.param sky130_fd_pr__nfet_01v8__u0_diff_60=0.0010868
.param sky130_fd_pr__nfet_01v8__nfactor_diff_60=0.32842233
.param sky130_fd_pr__nfet_01v8__keta_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_60=0.014447
.param sky130_fd_pr__nfet_01v8__ua_diff_60=2.61524e-11
.param sky130_fd_pr__nfet_01v8__ub_diff_60=1.86252e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_60=-2.39489e-11
.param sky130_fd_pr__nfet_01v8__tvoff_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_60=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_61=-26841.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_61=-0.037283
.param sky130_fd_pr__nfet_01v8__pdits_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__b1_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__voff_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__u0_diff_61=0.0035962
.param sky130_fd_pr__nfet_01v8__nfactor_diff_61=0.2721
.param sky130_fd_pr__nfet_01v8__keta_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_61=0.0062338
.param sky130_fd_pr__nfet_01v8__ua_diff_61=-3.67e-13
.param sky130_fd_pr__nfet_01v8__ub_diff_61=3.73839e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_61=0.0
.param sky130_fd_pr__nfet_01v8__tvoff_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__rdsw_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__a0_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__vsat_diff_62=-36357.0
.param sky130_fd_pr__nfet_01v8__kt1_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__vth0_diff_62=-0.025691
.param sky130_fd_pr__nfet_01v8__pdits_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__b0_diff_62=-7.73903e-17
.param sky130_fd_pr__nfet_01v8__b1_diff_62=2.98947e-18
.param sky130_fd_pr__nfet_01v8__voff_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pditsd_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__pclm_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__u0_diff_62=0.0020168
.param sky130_fd_pr__nfet_01v8__nfactor_diff_62=-0.0492
.param sky130_fd_pr__nfet_01v8__keta_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__ags_diff_62=0.0
.param sky130_fd_pr__nfet_01v8__k2_diff_62=-0.0016789
.param sky130_fd_pr__nfet_01v8__ua_diff_62=3.9629e-12
.param sky130_fd_pr__nfet_01v8__ub_diff_62=2.0374e-19
.param sky130_fd_pr__nfet_01v8__eta0_diff_62=0.0
.include "sky130_fd_pr__nfet_01v8__ff.pm3.spice"