* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.model sky130_fd_pr__diode_pd2nw_11v0 d level=3.0 tlevc=1.0 area=1.0e+12 cj='0.00077547*1e-12*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult' mj=0.33956 pb=0.6587 cjsw='9.8717e-011*1e-6*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult' mjsw=0.24676 php=1 cta=0.00096 ctp=3e-005 tpb=0.001671 tphp=0 js=2.1483e-017 jsw=4.02e-018 n=1.3632 rs=600 ik='4.76e-008/1e-12' ikr='0/1e-12' vb=12.69 ibv=0.00106 trs=0 eg=1.05 xti=10.0 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0