* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_b__toxe_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_b__overlap_mult=0.9642
.param sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult=9.9543e-1
.param sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult=1.0204
.param sky130_fd_pr__rf_nfet_01v8_b__lint_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_b__wint_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_b__rshg_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_b__dlc_diff=-.61492e-9
.param sky130_fd_pr__rf_nfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_b__xgw_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_0=-0.019045
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_0=876.33
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_0=0.0076402
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_0=0.00078682
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_1=-0.0024718
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_1=292.74
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_1=0.01684
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_1=0.00069507
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_2=-0.011464
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_2=4008.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_2=0.034561
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_2=-0.00018668
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_3=0.0031296
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_3=-7677.3
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_3=0.0045864
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_3=-0.0050888
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_4=-0.019118
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_4=-3226.1
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_4=0.020455
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_4=-0.0033825
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_5=-0.010928
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_5=-3103.8
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_5=0.037245
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_5=-0.00010837
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_6=-0.0038131
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_6=-0.010357
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_6=-10521.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_6=0.0019487
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_7=0.017771
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_7=-0.0036526
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_7=-0.018633
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_7=-3856.6
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_8=0.03546
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_8=-0.0023259
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_8=-0.014738
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_8=-749.49
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_0=0.0066076
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_0=-0.00069668
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_0=0.0055162
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_0=-9578.4
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_1=0.022438
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_1=-0.0013475
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_1=-0.017125
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_1=-1947.1
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_2=0.0375
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_2=-0.0010013
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_2=-0.013525
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_2=3934.3
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_3=-9286.3
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_3=0.0055484
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_3=-0.005738
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_3=-0.0050065
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_4=-2375.7
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_4=0.023623
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_4=-0.0067253
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_4=-0.025509
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_5=14291.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_5=0.039092
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_5=-0.0049774
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_5=-0.018429
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_6=-11321.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_6=0.0029951
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_6=-0.0037175
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_6=-0.011302
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_7=-0.0055361
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_7=-8608.4
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_7=0.021579
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_7=-0.029895
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_8=-0.019214
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_8=-0.0040927
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_8=9127.9
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_8=0.037329
.include "sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"