* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_05v0_nvt__toxe_mult=0.9635
.param sky130_fd_pr__nfet_05v0_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_05v0_nvt__overlap_mult=5.1025e-1
.param sky130_fd_pr__nfet_05v0_nvt__ajunction_mult=6.8772e-1
.param sky130_fd_pr__nfet_05v0_nvt__pjunction_mult=9.0190e-1
.param sky130_fd_pr__nfet_05v0_nvt__lint_diff=1.21275e-8
.param sky130_fd_pr__nfet_05v0_nvt__wint_diff=-2.252e-8
.param sky130_fd_pr__nfet_05v0_nvt__dlc_diff=1.6112e-8
.param sky130_fd_pr__nfet_05v0_nvt__dwc_diff=-2.252e-8
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0=0.056665
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_0=-0.052927
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_0=-0.00059672
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_0=-0.0090633
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_0=-3.141e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0=-0.030851
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_0=-0.005637
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_0=-1.5907e-18
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_1=-1.357e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1=-0.019967
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_1=-0.032965
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_1=-0.0051327
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_1=-0.0077525
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_1=-2.636e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1=-0.018137
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_1=-0.0051202
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_2=-1.8782e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2=0.066292
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_2=0.00087158
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_2=-0.0096682
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_2=-4.2384e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2=-6160.2
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2=-0.03046
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_3=-2.0373e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_3=-0.0020789
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_3=-1.0928e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3=0.015653
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_3=0.0012297
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_3=-0.0052343
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_3=-0.0065532
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3=-0.024011
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_4=-0.0083037
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4=-0.020154
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_4=-2.6021e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_4=-0.038115
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_4=-1.4421e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4=-0.05753
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_4=-0.17718
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_4=-0.0022264
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_5=-0.00093844
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_5=-0.007664
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5=-0.017363
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_5=-2.4895e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_5=-0.0093971
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_5=-1.3242e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5=-0.0035696
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_5=-0.044469
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_6=-0.047321
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_6=-0.0028201
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_6=-0.0068477
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6=-0.023509
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_6=-2.2313e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_6=-0.009358
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_6=-1.1832e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6=-0.022424
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7=0.043963
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_7=-3.5325e-6
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_7=-0.010425
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7=-0.038579
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_7=-3.6456e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7=-6428.9
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_7=-1.7165e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8=0.017354
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_8=1.5203e-7
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_8=-0.0095342
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_8=-0.0085304
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8=-0.055166
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_8=-3.4036e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_8=-4.5502e-9
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_8=-1.6434e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9=-0.13265
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_9=-0.0070168
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_9=-0.0087887
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9=-0.042098
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_9=-2.2834e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9=-8459.3
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_9=-1.3613e-18
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10=-7916.1
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10=-0.035797
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10=0.028686
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_10=-0.010001
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_10=0.00041829
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_10=-3.5554e-11
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_10=-1.6633e-18
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10=0.0
.include "sky130_fd_pr__nfet_05v0_nvt.pm3.spice"