* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_20v0_zvt__cjdnwpsubjunction_mult=7.0510e-1
.param sky130_fd_pr__nfet_20v0_zvt__mjdnwpsubjunction_mult=1.6541
.param sky130_fd_pr__nfet_20v0_zvt__pbdnwpsubjunction_mult=1.4206
.param sky130_fd_pr__nfet_20v0_zvt__vb=30.0
.param n20zvtvh1defet_js_mult='max(0.1,n20zvtvh1defet_js_mult_pmc)'
.model sky130_fd_pr__nfet_20v0_zvt__parasitic__diode_ps2dn__extended_drain d level=3.0 tlevc=1.0 scalm=1.0e-6 area=1.0e+12 cj='1.6920e-004*sky130_fd_pr__nfet_20v0_zvt__cjdnwpsubjunction_mult*1e-12*sky130_fd_pr__model__parasitic__diode_ps2dn__ajunction_mult' mj='0.56056*sky130_fd_pr__nfet_20v0_zvt__mjdnwpsubjunction_mult' pb='0.21294*sky130_fd_pr__nfet_20v0_zvt__pbdnwpsubjunction_mult' cjsw='8.1380e-010*sky130_fd_pr__nfet_20v0_zvt__cjdnwpsubjunction_mult*1e-6*sky130_fd_pr__model__parasitic__diode_ps2dn__pjunction_mult' mjsw='0.18742*sky130_fd_pr__nfet_20v0_zvt__mjdnwpsubjunction_mult' php='0.21294*sky130_fd_pr__nfet_20v0_zvt__pbdnwpsubjunction_mult' cta=0.0031223 ctp=0.0014703 tpb=0.0016859 tphp=0.0016859 js='6.1049e-017*n20zvtvh1defet_js_mult' jsw='8.1115e-016*n20zvtvh1defet_js_mult' n=0.9891 rs=900 ik='2.08e-009/1e-12' ikr='0/1e-12' vb='sky130_fd_pr__nfet_20v0_zvt__vb' ibv=0.00106 trs=0 eg=1.17 xti=1.0 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0