* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap c0 c1 b
.param mult=1.0
.param ctot_a='91.27e-15*sky130_fd_pr__model__cap_vpp_finger__cor+0.0283/sqrt(mult*2*41.1*2.7)*91.27e-15*sky130_fd_pr__model__cap_vpp_finger__cor*sky130_fd_pr__model__cap_vpp_only_p__slope'
.param c0_sub='4.434e-15*cli2s_vpp'
.param c1_sub='3.315e-15*cli2s_vpp'
.param rat_m4=0.125
.param rat_m3=0.125
.param rat_m2=0.375
.param rat_m1=0.375
.param cap_m4='rat_m4*ctot_a'
.param cap_m3='rat_m3*ctot_a'
.param cap_m2='rat_m2*ctot_a'
.param cap_m1='rat_m1*ctot_a'
.param lm1='41.1-0.96'
.param lm2='41.1-0.96'
.param lm3='41.1-0.96'
.param lm4='41.1-0.96'
.param wm1=0.160
.param wm2=0.160
.param wm3=0.300
.param wm4=0.300
.param nfm1=9.0
.param nfm2=9.0
.param nfm3=5.0
.param nfm4=5.0
.param nvia3=5.0
.param nvia2=5.0
.param nvia=5.0
ccmvpp_hd5_atlas_fingercap_l40 a2 a1 c='cap_m4'
rsm4 a0 a2 r='rm4*lm4/wm4*(1/3)*(1/nfm4)'
rvia3_0 a0 b0 r='rcvia3/nvia3'
rvia3_1 a1 b1 r='rcvia3/nvia3'
rsm3 b0 b2 r='rm3*lm3/wm3*(1/3)*(1/nfm3)'
cm3 b2 b1 c='cap_m3'
rvia2_0 b0 c0 r='rcvia2/nvia2'
rvia2_1 b1 c1 r='rcvia2/nvia2'
rsm2 c0 c2 r='(rm2*lm2/wm2*(1/3)*(1/nfm2)+rm2*lm2/wm2)'
cm2 c2 c1 c='cap_m2'
rvia_0 c0 d0 r='rcvia/nvia'
rvia_1 c1 d1 r='rcvia/nvia'
rsm1 d0 d2 r='rm1*lm1/wm1*(1/3)*(1/nfm1)'
cm1 d2 d1 c='cap_m1'
cm12b_0 d0 b c='c0_sub'
cm12b_1 d1 b c='c1_sub'
.ends sky130_fd_pr__cap_vpp_02p7x41p1_m1m2m3m4_shieldl1_fingercap