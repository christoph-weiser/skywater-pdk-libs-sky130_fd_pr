* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_lvt_b__toxe_mult=1.052
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rbpb_mult=1.2
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__overlap_mult=9.8026e-1
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__ajunction_mult=1.1755e+0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__pjunction_mult=1.0477e+0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__lint_diff=-1.7325e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__wint_diff=3.2175e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__rshg_diff=7.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dlc_diff=-1.5633e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_b__xgw_diff=6.4250e-8
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult_p42=1.15
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult_p42=1.35
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult_p42=1.35
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_cap_mult=1.15
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_dist_mult=1.35
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rgate_stub_mult=1.35
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rd_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt__aw_rs_mult=1.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_0=0.053368
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_0=-0.0019719
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_0=26569.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_0=-0.024863
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_1=-0.017808
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_1=0.047766
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_1=-0.00047355
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_1=30213.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_2=0.00040478
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_2=0.015345
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_2=-0.001204
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_2=18070.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_3=-0.029988
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_3=0.037878
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_3=-0.0051828
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_3=28757.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_4=-0.022408
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_4=0.020083
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_4=-0.0014964
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_4=25513.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_5=-0.0063582
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_5=0.012
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_5=-0.0026836
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_5=24731.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_6=-0.034961
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_6=0.032444
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_6=-0.0082913
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_6=19960.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_7=-0.021804
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_7=0.01554
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_7=-0.0040633
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_7=23539.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__k2_diff_8=-0.0057548
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vth0_diff_8=0.0080085
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__u0_diff_8=-0.0040879
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__vsat_diff_8=26010.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_0=-0.023869
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_0=0.050138
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_0=-0.0074552
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_0=34785.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_1=-0.017943
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_1=0.040645
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_1=-0.0035828
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_1=30760.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_2=-0.0065733
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_2=0.009983
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_2=-0.0036611
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_2=24896.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_3=-0.030893
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_3=0.041356
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_3=-0.0055014
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_3=28064.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_4=-0.0064683
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_4=30230.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_4=-0.022603
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_4=0.021578
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_5=-0.0014353
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_5=-0.0058089
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_5=37969.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_5=-0.0073485
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_6=-0.035237
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_6=0.031623
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_6=-0.0062253
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_6=24780.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_7=-0.02312
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_7=0.012306
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_7=-0.0086402
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_7=24437.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__pclm_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__k2_diff_8=-0.0069151
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__u0_diff_8=-0.0086411
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vsat_diff_8=52788.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__vth0_diff_8=-0.0097748
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_lvt_bm04__ua_diff_8=0.0
.include "sky130_fd_pr__rf_nfet_01v8_lvt_b.pm3.spice"