* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__esd_rf_diode_pw2nd_11v0_200__parasitic__diode_pw2dn c0 c1
.param area=-1
.param perim=-1.0
resd_ndiode_h_dnwl_200 c0 a1 r=5.82
d1 a1 c1 sky130_fd_pr__model__parasitic__diode_pw2dn_noresistor area='area*1.65'
.ends sky130_fd_pr__esd_rf_diode_pw2nd_11v0_200__parasitic__diode_pw2dn