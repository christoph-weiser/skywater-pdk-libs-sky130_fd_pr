* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre=0.0
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm02 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm02 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__model.0 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.8292+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_0' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_0' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.0868e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_0' ua='1.663e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_0' ub='1.238e-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_0' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_0' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.0636+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_0' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_0' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_0' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_0' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_0' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.627+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_0' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3307+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_0' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.604e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='200*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=200.0 rbps=200.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='9e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.7e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='4.1e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='8e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='3.948e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.1869 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm02
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm02w5p00 d g s b
.param l=1
.param w=5.05
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm02w5p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__model l='l' w=5.05 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__model.1 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=4.995e-06 wmax=5.095e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.815+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_1' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_1' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.035e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_1' ua='1.512e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_1' ub='8.845e-19+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_1' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_1' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.0626+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_1' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_1' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_1' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_1' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_1' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.7788+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_1' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_1' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.004e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='140*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=140.0 rbps=140.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.21e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='2.755e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='5e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='3.748e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.1569 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm02w5p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm04 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm04 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__model.0 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.8372+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_0' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_0' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.0868e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_0' ua='1.663e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_0' ub='1.238e-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_0' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_0' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.0636+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_0' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_0' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_0' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_0' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_0' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.627+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_0' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3307+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_0' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.604e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='400*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=400.0 rbps=400.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.25e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.6e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='3.7e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2.1e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='3.348e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.3069 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm04
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm04w5p00 d g s b
.param l=1
.param w=5.05
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm04w5p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__model l='l' w=5.05 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__model.1 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=4.995e-06 wmax=5.095e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.50e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.815+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_1' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_1' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.035e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_1' ua='1.512e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_1' ub='8.845e-19+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_1' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_1' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.06175+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_1' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_1' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_1' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_1' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_1' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.6181+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_1' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_1' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.004e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='280*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=280.0 rbps=280.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='9e-7+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.3e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='3.755e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1.00e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='3.348e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.3069 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm04w5p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm04w7p00 d g s b
.param l=1
.param w=7.09
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm04w7p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__model l='l' w=7.09 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__model.2 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=7.085e-06 wmax=7.095e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.811+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_2' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_2' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.056e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_2' ua='1.588e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_2' ub='8.757e-19+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_2' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_2' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.06298+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_2' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_2' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_2' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_2' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_2' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.7232+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_2' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_2' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.004e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='220*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=220.0 rbps=220.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.5e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.3e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='3.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='3.348e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.3069 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm04w7p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm10 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm10 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__model.0 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=3.005e-06 wmax=3.015e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.8292+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_0' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_0' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.0868e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_0' ua='1.663e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_0' ub='1.238e-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_0' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_0' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.06175+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_0' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_0' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_0' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_0' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_0' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.7376+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_0+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_0' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3307+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_0' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.604e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='1000*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=1000.0 rbps=1000.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.25e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.7e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='3.7e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2.2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='3.048e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.2969 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm10
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm10w5p00 d g s b
.param l=1
.param w=5.05
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm10w5p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__model l='l' w=5.05 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__model.1 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=5.045e-06 wmax=5.055e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.815+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_1' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_1' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.056e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_1' ua='1.724e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_1' ub='1.624e-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_1' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_1' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.06545+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_1' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_1' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_1' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_1' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_1' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.7664+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_1+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_1' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3207+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_1' kt2=-0.01915 at=4.0e+4 ute=-1.377 ua1=3.094e-9 ub1=-1.812e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='700*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=700.0 rbps=700.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.25e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.3e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='3.6e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='2e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='2.848e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.3069 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm10w5p00
.subckt sky130_fd_pr__rf_nfet_g5v0d10v5_bm10w7p00 d g s b
.param l=1
.param w=7.09
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__rf_nfet_g5v0d10v5_bm10w7p00 d g s b sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__model l='l' w=7.09 ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__model.2 nmos lmin=4.95e-07 lmax=5.05e-07 wmin=7.085e-06 wmax=7.095e-6 level=54.0 tnom=30.0 version=4.5 toxm=1.16e-8 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='7.345e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='2.135e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff' wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-4.129e-9 dwb=-1.694e-9 igcmod=0.0 igbmod=0.0 rgatemod=3.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=1.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.794 rnoib=0.38 tnoia=7.5e+6 tnoib=7.2e+6 epsrox=3.9 toxe='1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult+sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope_spectre*(1.16e-08*sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_toxe_slope1/sqrt(l*w*mult)))' dtox=0.0 ndep=6.0e+17 nsd=1.0e+20 rshg='49.2+sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff' rsh=1.0 vth0='0.811+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_2' k1=0.8833 k2='-0.03308+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_2' k3=-0.884 dvt0=0.0 dvt1=0.53 dvt2=-0.1925 dvt0w=0.16 dvt1w=6.909e+6 dvt2w=-0.03602 w0=0.0 k3b=0.43 phin=0.0 lpe0=2.5e-8 lpeb=-2.182e-7 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat='1.056e+05+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_2' ua='1.89e-09+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_2' ub='1.437e-18+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_2' uc=6.62e-11 rdsw='724.6+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_2' prwb=0.05626 prwg=0.048 wr=1.0 u0='0.0655+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_2' a0='0.1745+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_2' keta=-0.01066 a1=0.0 a2=0.6597 ags='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_2' b0='3.293e-08+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_2' b1='0+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_2' eu=1.67 rdswmin=0.0 rdw=370.0 rdwmin=0.0 rsw=370.0 rswmin=0.0 voff='-0.2309+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_voff_slope/sqrt(l*w*mult))' nfactor='0.687+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_2+sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope_spectre*(sky130_fd_pr__rf_nfet_g5v0d10v5__b_nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-0.0008 cdsc=0.0 cdscb=0.0 cdscd=0.0 eta0=0.05 etab=-0.01932 dsub=0.2822 voffl=-4.258e-7 minv=0.0 pclm='0.5653+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_2' pdiblc1=0.211 pdiblc2=0.015 pdiblcb=-0.2683 drout=0.3896 pscbe1=9.373e+8 pscbe2=1.68e-6 pvag=1.99 delta=0.03542 alpha0=1.447e-5 alpha1=0.0 beta0=36.96 fprout=10.13 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=5.06e-11 bgidl=1.058e+9 cgidl=4000.0 egidl=0.8 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=1.16e-8 kt1='-0.3507+sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_2' kt2=-0.01915 at=4.0e+4 ute=-1.299 ua1=3.004e-9 ub1=-3.553e-18 uc1=-5.982e-11 kt1l=0.0 prt=0.0 xrcrg1=10.0 xrcrg2=2.0 rbpb='550*sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult' rbpd=550.0 rbps=550.0 rbdb=1.0e+5 rbsb=1.0e+5 gbmin=1.0e-12 noia=2.6e+41 noib=0.0 noic=0.0 em=4.1e+7 af=1.0 ef=0.89 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw='1.5e-06+sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff' xgl=0.0 ngcon=2.0 diomod=1.0 njs=1.077 jss=0.000375 jsws=5.84e-11 xtis=0.76 bvs=12.64 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001344 tpbsw=0.0009901 tpbswg=0.0 tcj=0.0006743 tcjsw=0.0002493 tcjswg=0.0 cgdo='2.3e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgso='3.4e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgbo=0.0 capmod=2.0 xpart=0.0 cgsl='5e-11*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cgdl='1.8e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult' cf=0.0 clc=1.0e-11 cle=0.6 dlc='1e-07+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff+sky130_fd_pr__rf_nfet_g5v0d10v5__base__dlc_rotweak' dwc='0+sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff' vfbcv=-1.0 acde=0.4176 moin=15.0 noff=2.0 voffcv=-0.1204 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs='0.001*sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult' mjs=0.295 pbs=0.985 cjsws='4.864e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjsws=0.03759 pbsws=0.8907 cjswgs='2.748e-10*sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult' mjswgs=0.3069 pbswgs=0.99
.ends sky130_fd_pr__rf_nfet_g5v0d10v5_bm10w7p00