* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__rf_nfet_20v0_nvt_aup d psub s
x0 d a_n900_n1000# s psub sky130_fd_pr__nfet_20v0_nvt w=3e+07u l=1.5e+06u
x1 d a_n900_n1000# s psub sky130_fd_pr__nfet_20v0_nvt w=3e+07u l=1.5e+06u
.ends