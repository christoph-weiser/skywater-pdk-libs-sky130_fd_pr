* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre=0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre=0.0
.subckt sky130_fd_pr__nfet_01v8 d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__nfet_01v8__model.0 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.5190093+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.026724591 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.63331 eta0=0.08 etab=-0.07 u0=0.0318614 ua=-7.5866357e-10 ub=1.674192e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.334619 ags=0.4051693 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.1 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.5190093+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.54086565 k2=-0.026724591 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.63331 eta0=0.08 etab=-0.07 u0=0.0318614 ua=-7.5866357e-10 ub=1.674192e-18 uc=4.9242e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.334619 ags=0.4051693 a1=0.0 a2=0.42385546 b0=0.0 b1=2.1073424e-24 keta=-0.0087946 dwg=0.0 dwb=0.0 pclm=0.026316 pdiblc1=0.39 pdiblc2=0.0030734587 pdiblcb=-0.025 drout=0.56 pscbe1=754674160.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31303 kt2=-0.045313337 at=140000.0 ute=-1.8134 ua1=3.7602e-10 ub1=-6.3962e-19 uc1=1.5829713e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.2 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.194724788e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-3.694376992e-09 wvth0=-4.629762938e-08 pvth0=3.692761884e-13 k1=5.415457968e-01 lk1=-5.424943089e-09 wk1=-6.798494173e-08 pk1=5.422571412e-13 k2=-2.716644654e-02 lk2=3.524299843e-09 wk2=4.416623650e-08 pk2=-3.522759090e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.049994782e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.146551938e-09 wvoff=-2.690041279e-08 pvoff=2.145613508e-13 nfactor=2.636374809e+00 lnfactor=-2.444533584e-08 wnfactor=-3.063469433e-07 pnfactor=2.443464883e-12 eta0=0.08 etab=-0.07 u0=3.183773360e-02 lu0=1.887663852e-10 wu0=2.365604853e-09 pu0=-1.886838603e-14 ua=-7.582789781e-10 lua=-3.067557542e-18 wua=-3.844237946e-17 pua=3.066216468e-22 ub=1.672091096e-18 lub=1.675709387e-26 wub=2.099985257e-25 pub=-1.674976801e-30 uc=4.877008480e-11 luc=3.764059839e-18 wuc=4.717088911e-17 puc=-3.762414268e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.327488969e+00 la0=5.687009899e-08 wa0=7.126914150e-07 pa0=-5.684523652e-12 ags=4.061230713e-01 lags=-7.607409863e-09 wags=-9.533543630e-08 pags=7.604084055e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=1.950656262e-24 lb1=1.249749944e-30 wb1=1.566176377e-29 pb1=-1.249203578e-34 keta=-8.288058846e-03 lketa=-4.040241132e-09 wketa=-5.063197041e-08 pketa=4.038474820e-13 dwg=0.0 dwb=0.0 pclm=6.800573404e-02 lpclm=-3.325229885e-07 wpclm=-4.167150812e-06 ppclm=3.323776161e-11 pdiblc1=0.39 pdiblc2=3.074732157e-03 lpdiblc2=-1.015726833e-11 wpdiblc2=-1.272900534e-10 ppdiblc2=1.015282777e-15 pdiblcb=-0.025 drout=0.56 pscbe1=7.580442487e+08 lpscbe1=-2.688028581e+01 wpscbe1=-3.368615365e+02 ppscbe1=2.686853428e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.131868837e-01 lkt1=1.251326022e-09 wkt1=1.568151505e-08 pkt1=-1.250778967e-13 kt2=-4.539671736e-02 lkt2=6.650530936e-10 wkt2=8.334390809e-09 pkt2=-6.647623457e-14 at=140000.0 ute=-1.816359229e+00 lute=2.360321122e-08 wute=2.957935066e-07 pute=-2.359289237e-12 ua1=3.613755352e-10 lua1=1.168062433e-16 wua1=1.463806258e-15 pua1=-1.167551779e-20 ub1=-6.204482125e-19 lub1=-1.529167842e-25 wub1=-1.916340595e-24 pub1=1.528499321e-29 uc1=1.690988400e-11 luc1=-8.615590785e-18 wuc1=-1.079698769e-16 puc1=8.611824221e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.3 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.124282658e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.431437174e-08 wvth0=4.256783852e-08 pvth0=1.593500235e-14 k1=5.304574419e-01 lk1=3.866386370e-08 wk1=1.369158390e-07 pk1=-2.724562297e-13 k2=-2.007149225e-02 lk2=-2.468620333e-08 wk2=-7.809516520e-08 pk2=1.338520518e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.378281302e-01 ldsub=8.815836977e-08 wdsub=2.216217672e-06 pdsub=-8.811982869e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.094030449e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.536262827e-08 wvoff=5.578493138e-08 pvoff=-1.142068228e-13 nfactor=2.592450448e+00 lnfactor=1.502038973e-07 wnfactor=1.313313239e-08 pnfactor=1.173168653e-12 eta0=7.412445450e-02 leta0=2.336196799e-08 weta0=5.872976830e-07 peta0=-2.335175460e-12 etab=-6.486356790e-02 letab=-2.042315258e-08 wetab=-5.134186554e-07 petab=2.041422399e-12 u0=3.209879152e-02 lu0=-8.492353878e-10 wu0=7.707681347e-09 pu0=-4.010920869e-14 ua=-7.772766349e-10 lua=7.246970951e-17 wua=1.349633081e-15 pua=-5.212555164e-21 ub=1.715448650e-18 lub=-1.556384353e-25 wub=-1.333196930e-24 pub=4.460978208e-30 uc=5.877915793e-11 luc=-3.603337616e-17 wuc=-3.264462550e-16 puc=1.109311150e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.442796403e+00 la0=-4.016079406e-07 wa0=-1.342075208e-06 pa0=2.485507888e-12 ags=4.028351540e-01 lags=5.465796758e-09 wags=-1.033597319e-06 pags=4.491065254e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=4.502912266e-24 lb1=-8.898367034e-30 wb1=-3.132352754e-29 pb1=6.189955043e-35 keta=-1.640202815e-02 lketa=2.822200432e-08 wketa=8.756343093e-08 pketa=-1.456362283e-13 dwg=0.0 dwb=0.0 pclm=-6.131369147e-01 lpclm=2.375792818e-06 wpclm=8.540188246e-06 ppclm=-1.728834668e-11 pdiblc1=0.39 pdiblc2=3.181248537e-03 lpdiblc2=-4.336808822e-10 wpdiblc2=-1.246582526e-08 ppdiblc2=5.007497679e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.031489705e+08 lpscbe1=1.913908060e+02 wpscbe1=6.737230730e+02 ppscbe1=-1.331368419e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.112847401e-01 lkt1=-6.311855597e-09 wkt1=3.394151730e-08 pkt1=-1.976821490e-13 kt2=-4.403955904e-02 lkt2=-4.731192969e-09 wkt2=-1.656662876e-08 pkt2=3.253360577e-14 at=1.381479098e+05 lat=7.364162488e-03 wat=1.851280495e-01 pat=-7.360943023e-7 ute=-1.757935204e+00 lute=-2.086986568e-07 wute=-1.613263360e-06 pute=5.231380497e-12 ua1=6.225548039e-10 lua1=-9.216780498e-16 wua1=-5.190223011e-15 pua1=1.478180753e-20 ub1=-9.463016587e-19 lub1=1.142720834e-24 wub1=5.188563162e-24 pub1=-1.296507040e-29 uc1=-2.357426518e-13 luc1=5.955775258e-17 wuc1=1.710346184e-16 puc1=-2.481773957e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.4 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.265214792e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.535734467e-09 wvth0=-1.282118392e-07 pvth0=3.534188715e-13 k1=5.524870904e-01 lk1=-4.869717742e-09 wk1=-2.472758915e-07 pk1=4.867588799e-13 k2=-3.352973142e-02 lk2=1.909107599e-09 wk2=8.620493828e-08 pk2=-1.908272975e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=5.824396194e-01 wdsub=-2.242980920e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.029956789e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.700801503e-09 wvoff=1.346030157e-07 pvoff=-2.699620766e-13 nfactor=2.660003227e+00 lnfactor=1.671041853e-08 wnfactor=1.452042175e-06 pnfactor=-1.670311306e-12 eta0=8.609480828e-02 leta0=-2.930790459e-10 weta0=-6.092143748e-07 peta0=2.929509176e-14 etab=-7.518471959e-02 letab=-2.715316148e-11 wetab=5.182452938e-07 petab=2.714129066e-15 u0=3.138075868e-02 lu0=5.696951655e-10 wu0=1.622703524e-08 pu0=-5.694461062e-14 ua=-7.784147269e-10 lua=7.471873419e-17 wua=2.491281076e-15 pua=-7.468606865e-21 ub=1.671533075e-18 lub=-6.885528766e-26 wub=-2.558588474e-24 pub=6.882518551e-30 uc=3.956352106e-11 luc=1.939335609e-18 wuc=3.330022481e-16 puc=-1.938487771e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.148217881e+04 lvsat=-2.928986896e-03 wvsat=-1.481530827e-01 pvsat=2.927706402e-7 a0=1.229249642e+00 la0=2.038950021e-08 wa0=9.470215552e-07 pa0=-2.038058633e-12 ags=4.282285224e-01 lags=-4.471495281e-08 wags=-1.022704940e-06 pags=4.469540432e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.862460185e-03 lketa=9.370520639e-09 wketa=4.878426501e-07 pketa=-9.366424034e-13 dwg=0.0 dwb=0.0 pclm=5.768770306e-01 lpclm=2.416342047e-08 wpclm=1.013853514e-06 ppclm=-2.415285670e-12 pdiblc1=4.131572185e-01 lpdiblc1=-4.576181312e-08 wpdiblc1=-2.314709462e-06 ppdiblc1=4.574180697e-12 pdiblc2=2.903299932e-03 lpdiblc2=1.155833635e-10 wpdiblc2=1.872041904e-08 ppdiblc2=-1.155328327e-14 pdiblcb=-2.318864550e-02 lpdiblcb=-3.579482830e-09 wpdiblcb=-1.810562609e-07 ppdiblcb=3.577917952e-13 drout=5.380958797e-01 ldrout=4.328552063e-08 wdrout=2.189454424e-06 pdrout=-4.326659707e-12 pscbe1=7.606510411e+08 lpscbe1=7.775889417e+01 wpscbe1=3.933175629e+03 ppscbe1=-7.772489954e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.205658464e-07 lalpha0=-3.765840295e-13 walpha0=-1.904825348e-11 palpha0=3.764193945e-17 alpha1=8.524824670e-01 lalpha1=-4.905692338e-09 walpha1=-2.481381680e-07 palpha1=4.903547668e-13 beta0=1.406239407e+01 lbeta0=-3.999582106e-07 wbeta0=-2.023055887e-05 pbeta0=3.997833569e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.107339048e-01 lkt1=-7.400381177e-09 wkt1=-4.404168957e-07 pkt1=7.397145879e-13 kt2=-4.496893626e-02 lkt2=-2.894617183e-09 wkt2=-1.465179912e-07 pkt2=2.893351714e-13 at=1.381088459e+05 lat=7.441358137e-03 wat=1.890327353e-01 pat=-7.438104924e-7 ute=-1.803083395e+00 lute=-1.194796923e-07 wute=-5.009469552e-06 pute=1.194274582e-11 ua1=2.816514627e-10 lua1=-2.480066846e-16 wua1=-1.025466117e-14 pua1=2.478982610e-20 ub1=-4.339323422e-19 lub1=1.302093822e-25 wub1=5.213953787e-24 pub1=-1.301524572e-29 uc1=3.132149136e-11 luc1=-2.803633615e-18 wuc1=-9.636508894e-17 puc1=2.802407923e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.5 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.173374665e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.429110907e-09 wvth0=1.451912490e-07 pvth0=8.654027462e-14 k1=5.406566785e-01 lk1=6.678373256e-09 wk1=9.474366135e-07 pk1=-6.794430059e-13 k2=-2.740120282e-02 lk2=-4.073169797e-09 wk2=-3.944736425e-07 pk2=2.783803696e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.991414420e-01 ldsub=-3.091440504e-07 wdsub=-5.343647045e-06 pdsub=3.026671828e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.009256027e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.801256000e-10 wvoff=-4.674916482e-08 pvoff=-9.293768455e-14 nfactor=2.605596465e+00 lnfactor=6.981881780e-08 wnfactor=-8.349209003e-07 pnfactor=5.620756817e-13 eta0=2.018846564e-01 leta0=-1.133197182e-07 weta0=-4.615884383e-06 peta0=3.940349927e-12 etab=-1.463451305e-01 letab=6.943508571e-08 wetab=1.015844159e-06 petab=-4.830100369e-13 u0=3.352698870e-02 lu0=-1.525317221e-09 wu0=-3.802867750e-08 pu0=-3.983656204e-15 ua=-5.371888159e-10 lua=-1.607505616e-16 wua=-5.221570888e-15 pua=6.018559916e-23 ub=1.475966341e-18 lub=1.220444419e-25 wub=5.223075908e-24 pub=-7.134441927e-31 uc=1.095109860e-11 luc=2.986895122e-17 wuc=2.023582373e-16 puc=-6.632245490e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.943645684e+04 lvsat=-9.320840406e-04 wvsat=5.632967890e-02 pvsat=9.316765521e-8 a0=1.291158855e+00 la0=-4.004231074e-08 wa0=-4.167785480e-06 pa0=2.954688648e-12 ags=2.381856961e-01 lags=1.407926915e-07 wags=2.198736236e-06 pags=1.324975729e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=3.561401696e-03 lketa=-8.045862015e-10 wketa=-7.306170793e-07 pketa=2.527400029e-13 dwg=0.0 dwb=0.0 pclm=6.404786183e-01 lpclm=-3.792037900e-08 wpclm=-2.690702931e-06 ppclm=1.200865240e-12 pdiblc1=3.871350928e-01 lpdiblc1=-2.036067943e-08 wpdiblc1=2.863654728e-07 ppdiblc1=2.035177815e-12 pdiblc2=1.217587306e-03 lpdiblc2=1.761068143e-09 wpdiblc2=2.331725074e-08 ppdiblc2=-1.604041618e-14 pdiblcb=-2.862270899e-02 lpdiblcb=1.724902169e-09 wpdiblcb=3.621125218e-07 ppdiblcb=-1.724148077e-13 drout=5.994456506e-01 ldrout=-1.660019935e-08 wdrout=-3.942840578e-06 pdrout=1.659294207e-12 pscbe1=8.616614397e+08 lpscbe1=-2.084099226e+01 wpscbe1=-6.163448258e+03 ppscbe1=2.083188100e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.410386908e-08 lalpha0=-2.336172208e-13 walpha0=-4.408458775e-12 palpha0=2.335150880e-17 alpha1=8.450350661e-01 lalpha1=2.363983782e-09 walpha1=4.962763360e-07 palpha1=-2.362950295e-13 beta0=1.380708182e+01 lbeta0=-1.507387305e-07 wbeta0=5.289504551e-06 pbeta0=1.506728306e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.095566483e-01 lkt1=-8.549543620e-09 wkt1=2.833493486e-07 pkt1=3.322030121e-14 kt2=-4.861045418e-02 lkt2=6.599995580e-10 wkt2=2.187908274e-07 pkt2=-6.725591757e-14 at=1.706731833e+05 lat=-2.434586389e-02 wat=-6.806270065e-01 pat=1.050956893e-7 ute=-2.105517726e+00 lute=1.757373462e-07 wute=1.205657763e-05 pute=-4.716037219e-12 ua1=-3.629341746e-10 lua1=3.811965610e-16 wua1=2.502228661e-14 pua1=-9.645272601e-21 ub1=-9.356348756e-20 lub1=-2.020369101e-25 wub1=-1.133769218e-23 pub1=3.141411760e-30 uc1=1.727110250e-11 luc1=1.091145677e-17 wuc1=7.294628321e-16 puc1=-5.258795712e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.6 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.254411003e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.570679116e-09 wvth0=6.566827542e-07 pvth0=-1.569992447e-13 k1=5.733572999e-01 lk1=-8.891569812e-09 wk1=-2.346183834e-06 pk1=8.887682595e-13 k2=-4.124433183e-02 lk2=2.518042280e-09 wk2=7.188101962e-07 pk2=-2.516941442e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.608544335e-01 ldsub=-5.232627283e-09 wdsub=-8.540599614e-08 pdsub=5.230339683e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.000421031e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.594596381e-10 wvoff=-1.874716975e-07 pvoff=-2.593462075e-14 nfactor=2.753747772e+00 lnfactor=-7.213529842e-10 wnfactor=1.941378547e-07 pnfactor=7.210376231e-14 eta0=-3.611397891e-02 weta0=3.659797201e-6 etab=-5.538291750e-04 letab=1.859865862e-11 wetab=5.311487409e-09 petab=-1.859052765e-15 u0=2.991463485e-02 lu0=1.946544869e-10 wu0=-5.531066347e-09 pu0=-1.945693879e-14 ua=-9.104153604e-10 lua=1.695603236e-17 wua=-1.535549350e-15 pua=-1.694861952e-21 ub=1.754640735e-18 lub=-1.064246927e-26 wub=1.490474610e-24 pub=1.063781659e-30 uc=7.380749713e-11 luc=-5.924295007e-20 wuc=5.062814353e-17 puc=5.921705023e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.910068385e+04 lvsat=-7.722104313e-04 wvsat=8.989229878e-02 pvsat=7.718728363e-8 a0=1.207060381e+00 wa0=2.037770596e-6 ags=4.506321897e-01 lags=3.963926782e-08 wags=1.330306265e-05 pags=-3.962193833e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.079528043e-03 lketa=3.771231919e-10 wketa=-1.206320433e-07 pketa=-3.769583212e-14 dwg=0.0 dwb=0.0 pclm=5.524057554e-01 lpclm=4.014281679e-09 wpclm=6.741296190e-07 ppclm=-4.012526715e-13 pdiblc1=2.847083853e-01 lpdiblc1=2.840836336e-08 wpdiblc1=1.052455833e-05 ppdiblc1=-2.839594379e-12 pdiblc2=4.856343117e-03 lpdiblc2=2.852550623e-11 wpdiblc2=-4.383054714e-09 ppdiblc2=-2.851303545e-15 pdiblcb=-3.853174870e-02 lpdiblcb=6.442952699e-09 wpdiblcb=1.352583289e-06 ppdiblcb=-6.440135969e-13 drout=5.984950270e-01 ldrout=-1.614757321e-08 wdrout=-3.847819773e-06 pdrout=1.614051381e-12 pscbe1=8.340729560e+08 lpscbe1=-7.705121978e+00 wpscbe1=-3.405805999e+03 ppscbe1=7.701753453e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.438818033e-07 lalpha0=1.082416053e-13 walpha0=6.735871957e-11 palpha0=-1.081942843e-17 alpha1=0.85 beta0=1.351261868e+01 lbeta0=-1.053422766e-08 wbeta0=3.472294548e-05 pbeta0=1.052962231e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.285216740e-01 lkt1=4.803878418e-10 wkt1=4.539688434e-07 pkt1=-4.801778259e-14 kt2=-4.748635604e-02 lkt2=1.247759616e-10 wkt2=1.037317342e-07 pkt2=-1.247214120e-14 at=1.176801617e+05 lat=8.860214216e-04 wat=-2.738963741e-01 pat=-8.856340708e-8 ute=-1.698659221e+00 lute=-1.798263502e-08 wute=-1.623367921e-06 pute=1.797477337e-12 ua1=4.605278602e-10 lua1=-1.088335838e-17 wua1=2.480129244e-15 pua1=1.087860040e-21 ub1=-4.886624463e-19 lub1=-1.391607233e-26 wub1=-7.661404497e-24 pub1=1.390998850e-30 uc1=4.720982253e-11 luc1=-3.343445632e-18 wuc1=-1.076907545e-15 puc1=3.341983944e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.7 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.226971824e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.191177740e-09 wvth0=9.309545878e-07 pvth0=-2.190219800e-13 k1=5.548884107e-01 lk1=-4.715089080e-09 wk1=-5.001023353e-07 pk1=4.713027737e-13 k2=-3.619588693e-02 lk2=1.376407145e-09 wk2=2.141864145e-07 pk2=-1.375805407e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.111893909e-01 ldsub=5.998426783e-09 wdsub=4.878927004e-06 pdsub=-5.995804390e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.009850091e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.726846397e-10 wvoff=-9.322231484e-08 pvoff=-4.724779914e-14 nfactor=2.807399696e+00 lnfactor=-1.285398430e-08 wnfactor=-5.168708917e-06 pnfactor=1.284836480e-12 eta0=-1.126962478e-01 leta0=1.731800795e-08 weta0=1.131467606e-05 peta0=-1.731043687e-12 etab=-5.054282121e-03 letab=1.036313086e-09 wetab=4.551600312e-07 petab=-1.035860031e-13 u0=3.278461961e-02 lu0=-4.543523865e-10 wu0=-2.924040723e-07 pu0=4.541537528e-14 ua=-6.073824236e-10 lua=-5.157062385e-17 wua=-3.182559504e-14 pua=5.154807821e-21 ub=1.544202603e-18 lub=3.694516816e-26 wub=2.252508788e-23 pub=-3.692901647e-30 uc=7.384766442e-11 luc=-6.832622020e-20 wuc=4.661317063e-17 puc=6.829634934e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.743328342e+04 lvsat=-3.951511689e-04 wvsat=2.565594458e-01 pvsat=3.949784167e-8 a0=1.207060381e+00 wa0=2.037770596e-6 ags=8.312126992e-01 lags=-4.642368628e-08 wags=-2.473835008e-05 pags=4.640339077e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.632681265e-03 lketa=2.589933484e-11 wketa=-2.758794648e-07 pketa=-2.588801217e-15 dwg=0.0 dwb=0.0 pclm=5.492089963e-01 lpclm=4.737183991e-09 wpclm=9.936657716e-07 ppclm=-4.735112989e-13 pdiblc1=4.531641189e-01 lpdiblc1=-9.685542409e-09 wpdiblc1=-6.313650481e-06 ppdiblc1=9.681308084e-13 pdiblc2=6.031854250e-03 lpdiblc2=-2.372998792e-10 wpdiblc2=-1.218827769e-07 ppdiblc2=2.371961364e-14 pdiblcb=1.309104138e-02 lpdiblcb=-5.230818559e-09 wpdiblcb=-3.807438874e-06 ppdiblcb=5.228531750e-13 drout=4.798565019e-01 ldrout=1.068086830e-08 wdrout=8.010846098e-06 pdrout=-1.067619884e-12 pscbe1=7.993153719e+08 lpscbe1=1.548190656e-01 wpscbe1=6.843288191e+01 ppscbe1=-1.547513818e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.040459718e-07 lalpha0=9.923328974e-14 walpha0=6.337687796e-11 palpha0=-9.918990693e-18 alpha1=9.069090007e-01 lalpha1=-1.286917378e-08 walpha1=-5.688412120e-06 palpha1=1.286354763e-12 beta0=1.277748789e+01 lbeta0=1.557053069e-07 wbeta0=1.082038852e-04 pbeta0=-1.556372356e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.209694650e-01 lkt1=-1.227438479e-09 wkt1=-3.009218830e-07 pkt1=1.226901867e-13 kt2=-4.630223396e-02 lkt2=-1.429966677e-10 wkt2=-1.462870566e-08 pkt2=1.429341524e-14 at=1.232736586e+05 lat=-3.788696079e-04 wat=-8.330015340e-01 pat=3.787039736e-8 ute=-1.937606266e+00 lute=3.605189395e-08 wute=2.226089029e-05 pute=-3.603613278e-12 ua1=7.614258198e-11 lua1=7.603999089e-17 wua1=4.090185251e-14 pua1=-7.600674773e-21 ub1=-2.691863256e-19 lub1=-6.354752435e-26 wub1=-2.959942151e-23 pub1=6.351974265e-30 uc1=3.935986943e-11 luc1=-1.568288639e-18 wuc1=-2.922554192e-16 puc1=1.567603014e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.8 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.0e-06 wmax=0.0001 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.273127829e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.470516334e-09 wvth0=4.695963186e-07 pvth0=-1.469873453e-13 k1=5.297223808e-01 lk1=-7.857658419e-10 wk1=2.015400442e-06 pk1=7.854223208e-14 k2=-2.971925463e-02 lk2=3.651716839e-10 wk2=-4.331936701e-07 pk2=-3.650120381e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.268343873e-01 ldsub=3.555679632e-09 wdsub=3.315111336e-06 pdsub=-3.554125160e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=3.701734074e-03 lcdscd=2.651605064e-10 wcdscd=1.697523848e-07 pcdscd=-2.650445835e-14 cit=0.0 voff='-1.177707254e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.093539242e-09 wvoff=1.584615478e-06 pvoff=-3.092186808e-13 nfactor=2.181380466e+00 lnfactor=8.489015405e-08 wnfactor=5.740584569e-05 pnfactor=-8.485304178e-12 eta0=-1.127808870e-02 leta0=1.482982266e-09 weta0=1.177293955e-06 peta0=-1.482333935e-13 etab=-2.892433920e-03 letab=6.987707553e-10 wetab=2.390697228e-07 petab=-6.984652667e-14 u0=2.594768345e-02 lu0=6.131394777e-10 wu0=3.909906465e-07 pu0=-6.128714254e-14 ua=-1.451257292e-09 lua=8.018862258e-17 wua=5.252499926e-14 pua=-8.015356571e-21 ub=2.213250091e-18 lub=-6.751723050e-26 wub=-4.435041155e-23 pub=6.748771332e-30 uc=6.294653549e-11 luc=1.633732446e-18 wuc=1.136249488e-15 puc=-1.633018211e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.018808429e+04 lvsat=-8.252747573e-04 wvsat=-1.880020667e-02 pvsat=8.249139637e-8 a0=1.207060381e+00 wa0=2.037770596e-6 ags=5.338841762e-01 wags=4.981503615e-6 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.221854762e-02 lketa=-3.032159495e-09 wketa=-2.233609846e-06 pketa=3.030833895e-13 dwg=0.0 dwb=0.0 pclm=5.427722098e-01 lpclm=5.742198078e-09 wpclm=1.637063011e-06 ppclm=-5.739687704e-13 pdiblc1=3.948535541e-01 lpdiblc1=-5.811640668e-10 wpdiblc1=-4.851432247e-07 ppdiblc1=5.809099935e-14 pdiblc2=4.739215410e-03 lpdiblc2=-3.547242126e-11 wpdiblc2=7.324595465e-09 ppdiblc2=3.545691343e-15 pdiblcb=6.744804231e-03 lpdiblcb=-4.239942475e-09 wpdiblcb=-3.173092604e-06 ppdiblcb=4.238088857e-13 drout=4.915551465e-01 ldrout=8.854288734e-09 wdrout=6.841493081e-06 pdrout=-8.850417816e-13 pscbe1=7.986209646e+08 lpscbe1=2.632410390e-01 wpscbe1=1.378432507e+02 ppscbe1=-2.631259553e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.786292971e-08 lalpha0=-9.917985016e-16 walpha0=-7.859492192e-13 palpha0=9.913649071e-20 alpha1=7.172123318e-01 lalpha1=1.674930532e-08 walpha1=1.327296161e-05 palpha1=-1.674198286e-12 beta0=1.341620656e+01 lbeta0=5.597832913e-08 wbeta0=4.435994207e-05 pbeta0=-5.595385653e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.150847439e-01 lkt1=-2.146255297e-09 wkt1=-8.891367274e-07 pkt1=2.145316997e-13 kt2=-4.510229766e-02 lkt2=-3.303499223e-10 wkt2=-1.345698772e-07 pkt2=3.302054999e-14 at=1.198289709e+05 lat=1.589701562e-04 wat=-4.886833555e-01 pat=-1.589006576e-8 ute=-1.132927038e+00 lute=-8.958750189e-08 wute=-5.817185347e-05 pute=8.954833602e-12 ua1=1.362272965e-09 lua1=-1.247712625e-16 wua1=-8.765495871e-14 pua1=1.247167150e-20 ub1=-1.134148121e-18 lub1=7.150415049e-26 wub1=5.685894360e-23 pub1=-7.147289030e-30 uc1=3.786297182e-11 luc1=-1.334569033e-18 wuc1=-1.426310994e-16 puc1=1.333985586e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.9 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.188270027e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.822538042e-08 wvth0=1.268111480e-09 pvth0=-1.267808858e-13 k1=5.418171603e-01 lk1=-9.512831965e-08 wk1=-6.618973728e-09 pk1=6.617394176e-13 k2=-2.674260415e-02 lk2=1.800885350e-09 wk2=1.253045661e-10 pk2=-1.252746634e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.045334456e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.349789870e-08 wvoff=-5.113941489e-09 pvoff=5.112721098e-13 nfactor=2.682355773e+00 lnfactor=-4.903406830e-06 wnfactor=-3.411762250e-07 pnfactor=3.410948067e-11 eta0=0.08 etab=-0.07 u0=3.155893251e-02 lu0=3.023953140e-08 wu0=2.104049190e-09 pu0=-2.103547080e-13 ua=-7.362717244e-10 lua=-2.238650203e-15 wua=-1.557639926e-16 pua=1.557268211e-20 ub=1.621184695e-18 lub=5.299465505e-24 wub=3.687337596e-25 pub=-3.686457650e-29 uc=4.772038059e-11 luc=1.521256295e-16 wuc=1.058481374e-17 puc=-1.058228778e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.349496651e+00 la0=-1.487410044e-06 wa0=-1.034931348e-07 pa0=1.034684372e-11 ags=4.021842899e-01 lags=2.984297781e-07 wags=2.076457219e-08 pags=-2.075961693e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=8.033273090e-25 lb1=1.303703901e-28 wb1=9.071096705e-30 pb1=-9.068931979e-34 keta=-7.180997052e-03 lketa=-1.613217878e-07 wketa=-1.122467714e-08 pketa=1.122199848e-12 dwg=0.0 dwb=0.0 pclm=5.760603957e-02 lpclm=-3.128257252e-06 wpclm=-2.176623391e-07 ppclm=2.176103961e-11 pdiblc1=0.39 pdiblc2=3.147856669e-03 lpdiblc2=-7.438021498e-09 wpdiblc2=-5.175332547e-10 ppdiblc2=5.174097506e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.174573788e+08 lpscbe1=3.720789982e+03 wpscbe1=2.588904254e+02 ppscbe1=-2.588286437e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.200657108e-01 lkt1=7.034031752e-07 wkt1=4.894238807e-08 pkt1=-4.893070846e-12 kt2=-4.543472374e-02 lkt2=1.213577724e-08 wkt2=8.444003956e-10 pkt2=-8.441988879e-14 at=140000.0 ute=-1.856901360e+00 lute=4.349097908e-06 wute=3.026077292e-07 pute=-3.025355149e-11 ua1=3.036703693e-10 lua1=7.233236521e-15 wua1=5.032844339e-16 pua1=-5.031643301e-20 ub1=-5.518932882e-19 lub1=-8.770577673e-24 wub1=-6.102517464e-25 pub1=6.101061160e-29 uc1=1.657054426e-11 luc1=-7.406544670e-17 wuc1=-5.153431152e-18 puc1=5.152201337e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.10 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.197393603e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=-5.078505592e-9 k1=5.370550621e-01 wk1=2.650752369e-8 k2=-2.665245232e-02 wk2=-5.018170326e-10 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.082127306e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=2.048020293e-8 nfactor=2.436892544e+00 wnfactor=1.366335211e-6 eta0=0.08 etab=-0.07 u0=3.307271532e-02 wu0=-8.426250962e-9 ua=-8.483379519e-10 wua=6.238002890e-16 ub=1.886474514e-18 wub=-1.476697033e-24 uc=5.533574872e-11 wuc=-4.238983453e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.275037304e+00 wa0=4.144670811e-7 ags=4.171236044e-01 wags=-8.315751231e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=7.329634002e-24 wb1=-3.632773307e-29 keta=-1.525672240e-02 wketa=4.495234571e-8 dwg=0.0 dwb=0.0 pclm=-9.899367781e-02 wpclm=8.716894561e-7 pdiblc1=0.39 pdiblc2=2.775511312e-03 wpdiblc2=2.072606052e-9 pdiblcb=-0.025 drout=0.56 pscbe1=9.037191254e+08 wpscbe1=-1.036798810e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.848535368e-01 wkt1=-1.960034236e-7 kt2=-4.482720999e-02 wkt2=-3.381636551e-9 at=140000.0 ute=-1.639186688e+00 wute=-1.211876929e-6 ua1=6.657642457e-10 wua1=-2.015542681e-15 ub1=-9.909460496e-19 wub1=2.443923075e-24 uc1=1.286284790e-11 wuc1=2.063835029e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.11 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.148619652e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.890276705e-08 wvth0=-1.422559663e-08 pvth0=7.295844208e-14 k1=5.247112438e-01 lk1=9.845597383e-08 wk1=4.912095597e-08 pk1=-1.803678113e-13 k2=-1.921302920e-02 lk2=-5.933785053e-08 wk2=-1.115997735e-08 pk2=8.501093616e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.176438305e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.522373547e-08 wvoff=6.105726766e-08 pvoff=-3.236481868e-13 nfactor=2.199884560e+00 lnfactor=1.890407919e-06 wnfactor=2.730002323e-06 pnfactor=-1.087679434e-11 eta0=0.08 etab=-0.07 u0=3.447003714e-02 lu0=-1.114522883e-08 wu0=-1.594544082e-08 pu0=5.997408090e-14 ua=-8.875308152e-10 lua=3.126076079e-16 wua=8.606698490e-16 pua=-1.889303825e-21 ub=2.069398670e-18 lub=-1.459027940e-24 wub=-2.553784995e-24 pub=8.591000067e-30 uc=1.754519487e-10 luc=-9.580631468e-16 wuc=-8.340638805e-16 puc=6.314499858e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.649897199e+00 la0=-2.989933508e-06 wa0=-1.530071156e-06 pa0=1.550990144e-11 ags=5.315577429e-01 lags=-9.127422523e-07 wags=-9.678943846e-07 pags=7.056781617e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=1.461553941e-23 lb1=-5.811337240e-29 wb1=-7.243873489e-29 pb1=2.880262616e-34 keta=-2.849915097e-02 lketa=1.056234113e-07 wketa=8.996208595e-08 pketa=-3.590038095e-13 dwg=0.0 dwb=0.0 pclm=-1.019244331e+00 lpclm=7.340044362e-06 wpclm=3.396067243e-06 ppclm=-2.013478054e-11 pdiblc1=0.39 pdiblc2=2.814622145e-03 lpdiblc2=-3.119533207e-10 wpdiblc2=1.682108545e-09 ppdiblc2=3.114661224e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.004186824e+09 lpscbe1=-8.013440292e+02 wpscbe1=-2.049098704e+03 ppscbe1=8.074241626e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.596744755e-01 lkt1=-2.008316174e-07 wkt1=-3.565658870e-07 pkt1=1.280668045e-12 kt2=-3.215028598e-02 lkt2=-1.011128700e-07 wkt2=-8.381152135e-08 pkt2=6.415196996e-13 at=140000.0 ute=-1.119515970e+00 lute=-4.144964319e-06 wute=-4.551644711e-06 pute=2.663844204e-11 ua1=1.919486860e-09 lua1=-9.999862079e-15 wua1=-9.374855506e-15 pua1=5.869887996e-20 ub1=-2.193186578e-18 lub1=9.589233961e-24 wub1=9.024070989e-24 pub1=-5.248415466e-29 uc1=-2.774183419e-11 luc1=3.238684666e-16 wuc1=2.026400666e-16 puc1=-1.451670441e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.12 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.169068434e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.077205303e-08 wvth0=1.141358972e-08 pvth0=-2.898644975e-14 k1=5.755339035e-01 lk1=-1.036218331e-07 wk1=-1.766487394e-07 pk1=7.173232021e-13 k2=-4.335284486e-02 lk2=3.664533954e-08 wk2=8.385648891e-08 pk2=-2.927874559e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.872126539e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.977631701e-08 wvoff=-8.808335947e-08 pvoff=2.693552298e-13 nfactor=2.672677676e+00 lnfactor=1.051818902e-08 wnfactor=-5.449500866e-07 pnfactor=2.144861831e-12 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386683513e-01 letab=2.730347037e-07 wetab=-1.176909134e-11 petab=4.679550776e-17 u0=3.338360510e-02 lu0=-6.825427303e-09 wu0=-1.229844233e-09 pu0=1.462867558e-15 ua=-4.089115672e-10 lua=-1.590447614e-15 wua=-1.212818208e-15 pua=6.355166684e-21 ub=1.219303835e-18 lub=1.921064737e-24 wub=2.118126316e-24 pub=-9.985154686e-30 uc=-2.097160150e-10 luc=5.734170597e-16 wuc=1.541281884e-15 puc=-3.130197947e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=5.067133469e-01 la0=1.555520962e-06 wa0=5.169582504e-06 pa0=-1.112883267e-11 ags=1.121682116e-02 lags=1.156204019e-06 wags=1.690610240e-06 pags=-3.513794328e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.528191736e-05 lketa=-7.632325869e-09 wketa=-2.642739693e-08 pketa=1.037766034e-13 dwg=0.0 dwb=0.0 pclm=8.347779938e-01 lpclm=-3.180054735e-08 wpclm=-1.531916169e-06 ppclm=-5.404482921e-13 pdiblc1=0.39 pdiblc2=1.329904060e-03 lpdiblc2=5.591487706e-09 wpdiblc2=4.126490088e-10 ppdiblc2=8.162204988e-15 pdiblcb=-0.025 drout=0.56 pscbe1=8.052652765e+08 lpscbe1=-1.040490249e+01 wpscbe1=-3.662674833e+01 ppscbe1=7.237943593e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.046813117e-01 lkt1=-2.187831584e-08 wkt1=-1.199379323e-08 pkt1=-8.939746185e-14 kt2=-5.814765051e-02 lkt2=2.256187043e-09 wkt2=8.157323401e-08 pkt2=-1.607258004e-14 at=1.677727274e+05 lat=-1.104281413e-01 wat=-2.095053599e-02 pat=8.330218036e-8 ute=-2.533689068e+00 lute=1.477980245e-06 wute=3.783099279e-06 pute=-6.501633589e-12 ua1=-1.721514169e-09 lua1=4.477253188e-15 wua1=1.111578179e-14 pua1=-2.277468066e-20 ub1=1.239867144e-18 lub1=-4.061054535e-24 wub1=-1.001904353e-23 pub1=2.323385853e-29 uc1=6.727091944e-11 luc1=-5.391516357e-17 wuc1=-2.985607600e-16 puc1=5.411722084e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.13 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.143687095e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.578775095e-08 wvth0=-4.367374611e-08 pvth0=7.987361772e-14 k1=4.340894578e-01 lk1=1.758916280e-07 wk1=5.763314291e-07 pk1=-7.706680160e-13 k2=1.029185668e-02 lk2=-6.936388639e-08 wk2=-2.186303863e-07 pk2=3.049677476e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.133108041e+00 ldsub=-1.725380231e-06 wdsub=-6.073585748e-06 pdsub=1.200223145e-11 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.040740042e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-9.437217258e-09 wvoff=1.421041504e-07 pvoff=-1.855265952e-13 nfactor=2.605050780e+00 lnfactor=1.441581330e-07 wnfactor=1.834306898e-06 pnfactor=-2.556873549e-12 eta0=-6.411041806e-03 leta0=1.365715851e-08 weta0=3.428240498e-08 peta0=-6.774669465e-14 etab=-9.632053257e-04 letab=9.106073408e-10 wetab=1.939510043e-09 petab=-3.809197436e-15 u0=3.384188646e-02 lu0=-7.731053598e-09 wu0=-8.932636692e-10 pu0=7.977385883e-16 ua=-9.299748179e-10 lua=-5.607557664e-16 wua=3.545575809e-15 pua=-3.048067035e-21 ub=2.074615850e-18 lub=2.308518719e-25 wub=-5.362545924e-24 pub=4.797671032e-30 uc=7.461009665e-11 luc=1.154999470e-17 wuc=8.920838520e-17 puc=-2.607032319e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.043538777e+04 lvsat=1.177077746e-01 wvsat=2.765056110e-01 pvsat=-5.464126921e-7 a0=2.240715045e+00 la0=-1.871102217e-06 wa0=-6.089017016e-06 pa0=1.111969115e-11 ags=1.178946725e+00 lags=-1.151389082e-06 wags=-6.244912459e-06 pags=1.216787776e-11 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.144506780e-02 lketa=-1.093249755e-07 wketa=8.223904274e-08 pketa=-1.109630600e-13 dwg=0.0 dwb=0.0 pclm=1.096795738e+00 lpclm=-5.495832446e-07 wpclm=-2.602847633e-06 ppclm=1.575857928e-12 pdiblc1=-1.884416637e-01 lpdiblc1=1.143079395e-06 wpdiblc1=1.870182013e-06 ppdiblc1=-3.695734003e-12 pdiblc2=6.815002987e-03 lpdiblc2=-5.247813747e-09 wpdiblc2=-8.490490509e-09 ppdiblc2=2.575601950e-14 pdiblcb=-4.898724213e-02 lpdiblcb=4.740205271e-08 wpdiblcb=-1.593947540e-09 ppdiblcb=3.149857116e-15 drout=8.528408000e-01 ldrout=-5.786932471e-7 pscbe1=2.326916344e+09 lpscbe1=-3.017394357e+03 wpscbe1=-6.962207507e+03 ppscbe1=1.375826889e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.850882118e-07 lalpha0=-7.017025985e-13 walpha0=-2.019271745e-11 palpha0=3.990355590e-17 alpha1=8.168113760e-01 lalpha1=6.558523468e-8 beta0=1.182421474e+01 lbeta0=4.022988540e-06 wbeta0=-4.661152279e-06 pbeta0=9.211070820e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.599484662e-01 lkt1=8.733709777e-08 wkt1=-9.806652819e-08 pkt1=8.069396833e-14 kt2=-8.698809060e-02 lkt2=5.924881895e-08 wkt2=1.457790957e-07 pkt2=-1.429520948e-13 at=1.562147447e+05 lat=-8.758799562e-02 wat=6.308299700e-02 pat=-8.275950939e-8 ute=-2.561971268e+00 lute=1.533869719e-06 wute=2.695685041e-07 pute=4.415810628e-13 ua1=-8.561527015e-10 lua1=2.767181240e-15 wua1=-2.339774547e-15 pua1=3.815328618e-21 ub1=-3.464362798e-19 lub1=-9.263032314e-25 wub1=4.605306503e-24 pub1=-5.665846047e-30 uc1=1.177503932e-11 luc1=5.575224298e-17 wuc1=3.960554356e-17 puc1=-1.270903981e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.14 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.410704426e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.723227935e-09 wvth0=-1.990202568e-08 pvth0=5.666918563e-14 k1=7.174267341e-01 lk1=-1.006840875e-07 wk1=-2.822257427e-07 pk1=6.740054740e-14 k2=-1.063608615e-01 lk2=4.450503134e-08 wk2=1.547920100e-07 pk2=-5.954329653e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.707103633e+00 ldsub=1.047052631e-06 wdsub=1.278612866e-05 pdsub=-6.407414734e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.070483564e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.533844985e-09 wvoff=-4.157563511e-09 pvoff=-4.275527082e-14 nfactor=2.540704899e+00 lnfactor=2.069684633e-07 wnfactor=-3.835168691e-07 pnfactor=-3.919759284e-13 eta0=-4.518150604e-01 leta0=4.484320556e-07 weta0=-6.856480996e-08 peta0=3.264617435e-14 etab=2.383608940e-04 letab=-2.622847026e-10 wetab=-3.831943721e-09 petab=1.824526356e-15 u0=2.910477426e-02 lu0=-3.106987844e-09 wu0=-7.266506832e-09 pu0=7.018890676e-15 ua=-1.278540520e-09 lua=-2.205082364e-16 wua=-6.451937388e-17 pua=4.758768363e-22 ub=2.255126144e-18 lub=5.464927589e-26 wub=-1.969794008e-25 pub=-2.446244123e-31 uc=8.709476103e-11 luc=-6.367356515e-19 wuc=-3.273185511e-16 puc=1.458837056e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.852060170e+05 lvsat=-4.313076834e-02 wvsat=-6.794332083e-01 pvsat=3.867136032e-7 a0=-7.961271919e-01 la0=1.093268817e-06 wa0=1.035196488e-05 pa0=-4.928943148e-12 ags=-1.191493484e+00 lags=1.162482941e-06 wags=1.214398778e-05 pags=-5.782189765e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.110229117e-02 lketa=2.005927328e-08 wketa=-1.416725565e-07 pketa=1.076051128e-13 dwg=0.0 dwb=0.0 pclm=2.650604639e-01 lpclm=2.623034991e-07 wpclm=-7.918838127e-08 ppclm=-8.875767193e-13 pdiblc1=6.792427227e-01 lpdiblc1=2.961014293e-07 wpdiblc1=-1.745617576e-06 ppdiblc1=-1.662218555e-13 pdiblc2=-1.452074582e-03 lpdiblc2=2.821978283e-09 wpdiblc2=4.188817168e-08 ppdiblc2=-2.342040629e-14 pdiblcb=2.297448426e-02 lpdiblcb=-2.284237904e-08 wpdiblcb=3.187895080e-09 ppdiblcb=-1.517871612e-15 drout=1.020293091e+00 ldrout=-7.421494565e-07 wdrout=-6.870374051e-06 pdrout=6.706419445e-12 pscbe1=-1.461636461e+09 lpscbe1=6.807484247e+02 wpscbe1=9.998067113e+03 ppscbe1=-2.797265733e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.045363005e-05 lalpha0=1.963972049e-11 walpha0=1.383882472e-10 palpha0=-1.148930326e-16 alpha1=9.163772480e-01 lalpha1=-3.160459735e-8 beta0=1.569617265e+00 lbeta0=1.403287030e-05 wbeta0=9.041675896e-05 pbeta0=-8.359790114e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.686553668e-01 lkt1=-1.777383129e-09 wkt1=-1.171499994e-09 pkt1=-1.388875692e-14 kt2=-1.757666685e-02 lkt2=-8.506170576e-09 wkt2=2.911051178e-09 pkt2=-3.493453254e-15 at=7.989657716e+04 lat=-1.309108480e-02 wat=-4.915933551e-02 pat=2.680427210e-8 ute=-6.803264328e-01 lute=-3.028715436e-07 wute=2.142545094e-06 pute=-1.386698813e-12 ua1=2.582253735e-09 lua1=-5.891710656e-16 wua1=4.534728970e-15 pua1=-2.895121747e-21 ub1=-1.239485765e-18 lub1=-5.456547926e-26 wub1=-3.366333665e-24 pub1=2.115558900e-30 uc1=1.498316505e-10 luc1=-7.900978524e-17 wuc1=-1.926657220e-16 puc1=9.963794597e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.15 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.000559132e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.836187806e-08 wvth0=1.376410746e-07 pvth0=-1.834275596e-14 k1=2.822878334e-01 lk1=1.065012081e-07 wk1=-3.214225439e-07 pk1=8.606355554e-14 k2=5.208510788e-02 lk2=-3.093679874e-08 wk2=6.958429471e-08 pk2=-1.897283582e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.873282620e-01 ldsub=4.981820621e-08 wdsub=-9.651936128e-07 pdsub=1.400848462e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.031062123e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.410841694e-09 wvoff=-1.661568897e-07 pvoff=3.437844034e-14 nfactor=3.336221671e+00 lnfactor=-1.718057102e-07 wnfactor=-3.857714841e-06 pnfactor=1.262214797e-12 eta0=0.49 etab=-2.569930338e-04 letab=-2.642886484e-11 wetab=3.246611503e-09 petab=-1.545828615e-15 u0=2.615389718e-02 lu0=-1.701969034e-09 wu0=2.062968544e-08 pu0=-6.263490727e-15 ua=-1.349419498e-09 lua=-1.867602034e-16 wua=1.518287228e-15 pua=-2.777543679e-22 ub=1.999102462e-18 lub=1.765513675e-25 wub=-2.100701032e-25 pub=-2.383914576e-31 uc=4.031218941e-12 luc=3.891280702e-17 wuc=5.360116115e-16 puc=-2.651788647e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.892861902e+04 lvsat=2.175580681e-02 wvsat=2.997776903e-01 pvsat=-7.952395719e-8 a0=1.5 ags=2.363013912e+00 lags=-5.299459918e-07 wags=-3.898278820e-12 pags=1.856110885e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.540973132e-02 lketa=-6.457959399e-09 wketa=6.363471476e-08 pketa=9.850929874e-15 dwg=0.0 dwb=0.0 pclm=1.211362672e+00 lpclm=-1.882650489e-07 wpclm=-3.909760516e-06 ppclm=9.362965747e-13 pdiblc1=3.226103049e+00 lpdiblc1=-9.165504588e-07 wpdiblc1=-9.936612421e-06 ppdiblc1=3.733805666e-12 pdiblc2=6.207590322e-03 lpdiblc2=-8.250639262e-10 wpdiblc2=-1.378271132e-08 ppdiblc2=3.086505259e-15 pdiblcb=6.042263145e-01 lpdiblcb=-2.995973005e-07 wpdiblcb=-3.118623057e-06 ppdiblcb=1.484888708e-12 drout=-1.929948742e+00 ldrout=6.625668886e-07 wdrout=1.374074810e-05 pdrout=-3.107277813e-12 pscbe1=-7.843924541e+08 lpscbe1=3.582881720e+02 wpscbe1=7.852695801e+03 ppscbe1=-1.775777218e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=4.138540030e-05 lalpha0=-9.804068065e-12 walpha0=-2.250088190e-10 palpha0=5.813339291e-17 alpha1=0.85 beta0=4.244059302e+01 lbeta0=-5.427272610e-06 wbeta0=-1.665082017e-04 pbeta0=3.873332194e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.143827816e-01 lkt1=-2.761851474e-08 wkt1=-3.400134792e-07 pkt1=1.474461077e-13 kt2=-1.068137071e-03 lkt2=-1.636647591e-08 wkt2=-2.191664868e-07 pkt2=1.022456574e-13 at=7.917893229e+04 lat=-1.274938825e-02 wat=-6.070965093e-03 pat=6.288347764e-9 ute=-1.212504931e+00 lute=-4.948220236e-08 wute=-5.005194258e-06 pute=2.016597211e-12 ua1=1.746611269e-09 lua1=-1.912916045e-16 wua1=-6.466229626e-15 pua1=2.342830675e-21 ub1=-2.103656553e-18 lub1=3.568973429e-25 wub1=3.572949936e-24 pub1=-1.188483836e-30 uc1=-1.358491248e-10 luc1=5.701311637e-17 wuc1=1.965021153e-16 puc1=-8.565887140e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.16 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.860493656e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.519449341e-08 wvth0=4.902589364e-07 pvth0=-9.808234876e-14 k1=4.580806325e-01 lk1=6.674812771e-08 wk1=1.733198696e-07 pk1=-2.581551488e-14 k2=1.599447514e-02 lk2=-2.277540741e-08 wk2=-1.488644617e-07 pk2=3.042629217e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.052696561e+00 ldsub=-1.006455195e-07 wdsub=-9.748341775e-07 pdsub=1.422649249e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.072898457e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.799385846e-08 wvoff=-3.732545739e-07 pvoff=8.121068225e-14 nfactor=2.261485732e+00 lnfactor=7.123077612e-08 wnfactor=-1.371177436e-06 pnfactor=6.999191745e-13 eta0=1.550355063e+00 leta0=-2.397844526e-07 weta0=-2.539778355e-07 peta0=5.743353180e-14 etab=7.951944849e-02 letab=-1.806675425e-08 wetab=-1.331586887e-07 petab=2.930032036e-14 u0=-1.379440254e-02 lu0=7.331779670e-09 wu0=3.161274110e-08 pu0=-8.747155001e-15 ua=-5.194822301e-09 lua=6.828238050e-16 wua=8.593040434e-17 pua=4.615307479e-23 ub=4.384694130e-18 lub=-3.629167898e-25 wub=2.765827803e-24 pub=-9.113491065e-31 uc=3.482642912e-10 luc=-3.893068301e-17 wuc=-1.862306271e-15 puc=2.771671479e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.842631280e+04 lvsat=1.734667633e-02 wvsat=3.192144735e-01 pvsat=-8.391931360e-8 a0=1.5 ags=-2.725049684e+00 lags=6.206483575e-07 wags=1.392242436e-11 pags=-2.173791649e-18 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.132303484e-01 lketa=1.340144366e-08 wketa=5.300964428e-07 pketa=-9.563285946e-14 dwg=0.0 dwb=0.0 pclm=1.175664524e+00 lpclm=-1.801924126e-07 wpclm=-3.364135541e-06 ppclm=8.129111254e-13 pdiblc1=-3.504829723e+00 lpdiblc1=6.055557544e-07 wpdiblc1=2.121927084e-05 ppdiblc1=-3.311661150e-12 pdiblc2=-8.867346784e-03 lpdiblc2=2.583922051e-09 wpdiblc2=-1.823973298e-08 ppdiblc2=4.094398308e-15 pdiblcb=-2.245021456e+00 lpdiblcb=3.447201932e-07 wpdiblcb=1.190062844e-05 ppdiblcb=-1.911504749e-12 drout=2.107148649e+00 ldrout=-2.503661669e-07 wdrout=-3.309056973e-06 pdrout=7.482969076e-13 pscbe1=8.184696982e+08 lpscbe1=-4.176663670e+00 wpscbe1=-6.481001347e+01 ppscbe1=1.465587721e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.095849207e-06 lalpha0=-1.145422138e-12 walpha0=3.763936372e-11 palpha0=-1.260816547e-18 alpha1=-2.783651019e+00 lalpha1=8.216993069e-07 walpha1=1.998416412e-05 palpha1=-4.519138937e-12 beta0=4.486413993e+01 lbeta0=-5.975323815e-06 wbeta0=-1.149999148e-04 pbeta0=2.708544396e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-5.848447432e-01 lkt1=5.615627142e-08 wkt1=1.534668965e-06 pkt1=-2.764870815e-13 kt2=-1.553590431e-01 lkt2=1.852425241e-08 wkt2=7.440012128e-07 pkt2=-1.155612335e-13 at=3.846530241e+04 lat=-3.542570839e-03 wat=-2.430506920e-01 pat=5.987799529e-8 ute=-6.059333123e-01 lute=-1.866498818e-07 wute=1.299739770e-05 pute=-2.054436924e-12 ua1=4.223758656e-09 lua1=-7.514638060e-16 wua1=1.204986547e-14 pua1=-1.844325005e-21 ub1=-4.489634735e-18 lub1=8.964529052e-25 wub1=-2.407922044e-25 pub1=-3.260594437e-31 uc1=-9.851794355e-11 luc1=4.857119238e-17 wuc1=6.668615295e-16 puc1=-1.920240679e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.17 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.976807890e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.396977344e-09 wvth0=6.757248246e-07 pvth0=-1.270402507e-13 k1=8.024594106e-01 lk1=1.297820280e-08 wk1=1.181647507e-07 pk1=-1.720381524e-14 k2=-2.242879796e-02 lk2=-1.677615125e-08 wk2=-4.839081427e-07 pk2=8.273867234e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.439592925e+00 ldsub=-1.610539701e-07 wdsub=-5.121179048e-06 pdsub=7.896586276e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=6.411402419e-02 lcdscd=-9.167371879e-09 wcdscd=-2.504924994e-07 pcdscd=3.911089689e-14 cit=0.0 voff='5.546602005e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.140782643e-07 wvoff=-3.093003668e-06 pvoff=5.058614268e-13 nfactor=2.804112867e+01 lnfactor=-3.953899554e-06 wnfactor=-1.224818553e-04 pnfactor=1.960965597e-11 eta0=7.206115648e-02 leta0=-8.969555154e-09 weta0=5.975626641e-07 peta0=-7.552259564e-14 etab=3.506506218e-02 letab=-1.112582418e-08 wetab=-2.497332410e-08 petab=1.240869027e-14 u0=6.862122419e-02 lu0=-5.536266624e-09 wu0=9.414146325e-08 pu0=-1.851013956e-14 ua=6.033562110e-09 lua=-1.070331223e-15 wua=4.584847861e-16 pua=-1.201607616e-23 ub=-5.149634739e-18 lub=1.125735182e-24 wub=6.867891660e-24 pub=-1.551828949e-30 uc=1.721098632e-10 luc=-1.142663524e-17 wuc=3.768785961e-16 puc=-7.245022046e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.279489769e+05 lvsat=-7.560554356e-03 wvsat=-1.046666644e+00 pvsat=1.293439006e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.086656882e+00 lketa=1.653883689e-07 wketa=5.480040346e-06 pketa=-8.684973007e-13 dwg=0.0 dwb=0.0 pclm=-8.711599916e-01 lpclm=1.393905800e-07 wpclm=1.147277413e-05 ppclm=-1.503664604e-12 pdiblc1=-1.280695971e-01 lpdiblc1=7.832193538e-08 wpdiblc1=3.152457680e-06 ppdiblc1=-4.907812111e-13 pdiblc2=-6.906294732e-03 lpdiblc2=2.277731228e-09 wpdiblc2=8.833404804e-08 ppdiblc2=-1.254560557e-14 pdiblcb=-5.667230242e-01 lpdiblcb=8.267738936e-08 wpdiblcb=8.161113285e-07 ppdiblcb=-1.808125852e-13 drout=-2.487432580e-01 ldrout=1.174733719e-07 wdrout=1.199121755e-05 pdrout=-1.640626755e-12 pscbe1=8.143741681e+08 lpscbe1=-3.537203979e+00 wpscbe1=2.825952501e+01 ppscbe1=1.243717468e-7 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.219442353e-05 lalpha0=2.803299886e-12 walpha0=1.538681049e-10 palpha0=-1.940830728e-17 alpha1=9.328519045e+00 lalpha1=-1.069446478e-06 walpha1=-4.662971627e-05 palpha1=5.881685892e-12 beta0=-2.395538075e+01 lbeta0=4.769880867e-06 wbeta0=3.043272422e-04 pbeta0=-3.838662102e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-5.269357921e-01 lkt1=4.711459942e-08 wkt1=5.845589058e-07 pkt1=-1.281406973e-13 kt2=-6.472487730e-02 lkt2=4.372996302e-09 wkt2=1.930320397e-09 pkt2=3.027473130e-16 at=2.162270652e+05 lat=-3.129758143e-02 wat=-1.159255683e+00 pat=2.029305778e-7 ute=-9.375262849e+00 lute=1.182558155e-06 wute=-8.358412305e-07 pute=1.054296695e-13 ua1=-1.321109607e-08 lua1=1.970744671e-15 wua1=1.372150595e-14 pua1=-2.105328263e-21 ub1=8.031610843e-18 lub1=-1.058564294e-24 wub1=-6.900660490e-24 pub1=7.137857510e-31 uc1=2.439604408e-10 luc1=-4.902012639e-18 wuc1=-1.576303213e-15 puc1=1.582147024e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.18 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.201595472e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.149972668e-07 wvth0=-5.336354696e-09 pvth0=5.335081228e-13 k1=5.438271891e-01 lk1=-2.960832397e-07 wk1=-1.658124366e-08 pk1=1.657728671e-12 k2=-2.786182868e-02 lk2=1.136966286e-07 wk2=5.672496930e-09 pk2=-5.671143245e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.061807979e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=9.119802101e-08 wvoff=3.050801169e-09 pvoff=-3.050073126e-13 nfactor=2.614138722e+00 lnfactor=1.916670325e-06 wnfactor=-3.073283702e-09 pnfactor=3.072550294e-13 eta0=0.08 etab=-0.07 u0=3.178890457e-02 lu0=7.247812509e-09 wu0=9.642427617e-10 pu0=-9.640126548e-14 ua=-7.611659229e-10 lua=2.501755769e-16 wua=-3.238132445e-17 pua=3.237359697e-21 ub=1.678526098e-18 lub=-4.333064184e-25 wub=8.453359517e-26 pub=-8.451342208e-30 uc=5.878403900e-11 luc=-9.539761888e-16 wuc=-4.424979731e-17 puc=4.423923754e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.352085454e+00 la0=-1.746228537e-06 wa0=-1.163239711e-07 pa0=1.162962115e-11 ags=4.118255806e-01 lags=-6.654692147e-07 wags=-2.702038349e-08 pags=2.701393534e-12 a1=0.0 a2=0.42385546 b0=7.777924617e-25 lb0=-7.776068493e-29 wb0=-3.854958778e-30 pb0=3.854038830e-34 b1=2.633549380e-24 lb1=-5.260814057e-29 keta=-9.250464793e-03 lketa=4.557560051e-08 wketa=-9.678114294e-10 pketa=9.675804709e-14 dwg=0.0 dwb=0.0 pclm=1.614369198e-02 lpclm=1.016988051e-06 wpclm=-1.216325199e-08 ppclm=1.216034935e-12 pdiblc1=0.39 pdiblc2=2.773573112e-03 lpdiblc2=2.998140236e-08 wpdiblc2=1.337521605e-09 ppdiblc2=-1.337202419e-13 pdiblcb=-9.427960644e-01 lpdiblcb=9.175770416e-05 wpdiblcb=4.548856114e-06 ppdiblcb=-4.547770575e-10 drout=0.56 pscbe1=8.062271626e+08 lpscbe1=-5.154069996e+03 wpscbe1=-1.810776562e+02 ppscbe1=1.810344439e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.072159914e-01 lkt1=-5.812621098e-07 wkt1=-1.474444443e-08 pkt1=1.474092582e-12 kt2=-4.362268116e-02 lkt2=-1.690252377e-07 wkt2=-8.136593605e-09 pkt2=8.134651888e-13 at=140000.0 ute=-1.761372561e+00 lute=-5.201502322e-06 wute=-1.708599392e-07 pute=1.708191652e-11 ua1=4.317087131e-10 lua1=-5.567542354e-15 wua1=-1.313097049e-16 pua1=1.312783691e-20 ub1=-6.481907438e-19 lub1=8.568698527e-25 wub1=-1.329744002e-25 pub1=1.329426672e-29 uc1=1.484440068e-11 luc1=9.850771891e-17 wuc1=3.401823218e-18 puc1=-3.401011407e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.19 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.144028149e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.137091856e-8 k1=5.290053417e-01 wk1=6.640420812e-8 k2=-2.217020600e-02 wk2=-2.271709376e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016154495e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.221778293e-8 nfactor=2.710086723e+00 wnfactor=1.230782050e-8 eta0=0.08 etab=-0.07 u0=3.215172812e-02 wu0=-3.861578682e-9 ua=-7.486422008e-10 wua=1.296800320e-16 ub=1.656834896e-18 wub=-3.385383246e-25 uc=1.102824735e-11 wuc=1.772106370e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.264669722e+00 wa0=4.658517386e-7 ags=3.785123705e-01 wags=1.082106509e-7 a1=0.0 a2=0.42385546 b0=-3.114886529e-24 wb0=1.543825604e-29 b1=0.0 keta=-6.968962479e-03 wketa=3.875870406e-9 dwg=0.0 dwb=0.0 pclm=6.705384049e-02 wpclm=4.871113007e-8 pdiblc1=0.39 pdiblc2=4.274434057e-03 wpdiblc2=-5.356477769e-9 pdiblcb=3.650569948e+00 wpdiblcb=-1.821716117e-5 drout=0.56 pscbe1=5.482158036e+08 wpscbe1=7.251759048e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.363138165e-01 wkt1=5.904823407e-8 kt2=-5.208403914e-02 wkt2=3.258525515e-8 at=140000.0 ute=-2.021758369e+00 wute=6.842562112e-7 ua1=1.529990390e-10 wua1=5.258662831e-16 ub1=-6.052960693e-19 wub1=5.325330192e-25 uc1=1.977567061e-11 wuc1=-1.362354849e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.20 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.094048492e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.986445368e-08 wvth0=1.282140888e-08 pvth0=6.819205193e-14 k1=5.143584298e-01 lk1=1.168257617e-07 wk1=1.004324218e-07 pk1=-2.714136603e-13 k2=-1.480876321e-02 lk2=-5.871586889e-08 wk2=-3.298876161e-08 pk2=8.192821975e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016965986e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.472565646e-10 wvoff=-1.798171089e-08 pvoff=4.597387324e-14 nfactor=2.903642792e+00 lnfactor=-1.543829529e-06 wnfactor=-7.580219357e-07 pnfactor=6.144254900e-12 eta0=0.08 etab=-0.07 u0=3.163537691e-02 lu0=4.118487520e-09 wu0=-1.896065341e-09 pu0=-1.567720172e-14 ua=-6.610039312e-10 lua=-6.990147567e-16 wua=-2.620612688e-16 pua=3.124581892e-21 ub=1.468911821e-18 lub=1.498900005e-24 wub=4.223971663e-25 pub=-6.069324963e-30 uc=-1.023161189e-10 luc=9.040500801e-16 wuc=5.426329932e-16 puc=-2.914658410e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.014825383e+00 la0=1.992792425e-06 wa0=1.617523854e-06 pa0=-9.185893417e-12 ags=2.290185375e-01 lags=1.192383143e-06 wags=5.315752334e-07 pags=-3.376813488e-12 a1=0.0 a2=0.42385546 b0=-6.211189646e-24 lb0=2.469653475e-29 wb0=3.078440744e-29 pb0=-1.224029907e-34 b1=0.0 keta=-9.975873028e-03 lketa=2.398352748e-08 wketa=-1.844503110e-09 pketa=4.562647714e-14 dwg=0.0 dwb=0.0 pclm=-3.557238492e-01 lpclm=3.372132351e-06 wpclm=1.074726238e-07 ppclm=-4.686896653e-13 pdiblc1=0.39 pdiblc2=5.687552554e-03 lpdiblc2=-1.127122532e-08 wpdiblc2=-1.255694473e-08 ppdiblc2=5.743190375e-14 pdiblcb=7.304211445e+00 lpdiblcb=-2.914194148e-05 wpdiblcb=-3.632563876e-05 ppdiblcb=1.444356800e-10 drout=0.56 pscbe1=3.005663900e+08 lpscbe1=1.975285403e+03 wpscbe1=1.438242589e+03 ppscbe1=-5.687516851e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.574596798e-01 lkt1=1.686622815e-07 wkt1=1.280851606e-07 pkt1=-5.506479151e-13 kt2=-6.250017945e-02 lkt2=8.308055170e-08 wkt2=6.661110936e-08 pkt2=-2.713948407e-13 at=140000.0 ute=-2.363712447e+00 lute=2.727472228e-06 wute=1.614943892e-06 pute=-7.423291513e-12 ua1=-4.847675260e-10 lua1=5.086912859e-15 wua1=2.541307231e-15 pua1=-1.607543110e-20 ub1=-1.851937603e-19 lub1=-3.350793150e-24 wub1=-9.281076705e-25 pub1=1.165026879e-29 uc1=2.776052890e-11 luc1=-6.368831567e-17 wuc1=-7.244529657e-17 puc1=4.691702624e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.21 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.091809945e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.075453062e-08 wvth0=4.970507577e-08 pvth0=-7.846242378e-14 k1=5.393348269e-01 lk1=1.751620993e-08 wk1=2.764092559e-09 pk1=1.169288997e-13 k2=-2.493727473e-02 lk2=-1.844352959e-08 wk2=-7.416269826e-09 pk2=-1.975148544e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.294571546e+00 ldsub=-2.920756371e-06 wdsub=-2.171600641e-06 pdsub=8.634579485e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.065550189e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.996499625e-08 wvoff=3.057518639e-10 pvoff=-2.673956575e-14 nfactor=2.291134361e+00 lnfactor=8.915872952e-07 wnfactor=1.346086179e-06 pnfactor=-2.221965121e-12 eta0=2.746614598e-01 leta0=-7.740004382e-07 weta0=-5.754741697e-07 peta0=2.288163563e-12 etab=-2.401757413e-01 letab=6.766418914e-07 wetab=5.030874809e-07 petab=-2.000344244e-12 u0=3.487846788e-02 lu0=-8.776483274e-09 wu0=-8.638805747e-09 pu0=1.113285115e-14 ua=-8.425297392e-10 lua=2.275654349e-17 wua=9.363157329e-16 pua=-1.640328046e-21 ub=2.041556609e-18 lub=-7.780135537e-25 wub=-1.957190308e-24 pub=3.392238460e-30 uc=1.663509328e-10 luc=-1.642066562e-16 wuc=-3.226119606e-16 puc=5.256731990e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.316192760e+00 la0=-3.181621248e-06 wa0=-3.798707738e-06 pa0=1.234978000e-11 ags=5.898905223e-01 lags=-2.424929469e-07 wags=-1.177459808e-06 pags=3.418542267e-12 a1=0.0 a2=0.42385546 b0=3.077719703e-24 lb0=-1.223743211e-29 wb0=-1.525404677e-29 pb0=6.065216449e-35 b1=0.0 keta=-1.066629930e-02 lketa=2.672875624e-08 wketa=2.636204881e-08 pketa=-6.652660941e-14 dwg=0.0 dwb=0.0 pclm=6.023645232e-01 lpclm=-4.373573176e-07 wpclm=-3.800094678e-07 ppclm=1.469605428e-12 pdiblc1=0.39 pdiblc2=3.244423889e-04 lpdiblc2=1.005323008e-08 wpdiblc2=5.396000590e-09 ppdiblc2=-1.395144844e-14 pdiblcb=-0.025 drout=0.56 pscbe1=7.825561225e+08 lpscbe1=5.882867629e+01 wpscbe1=7.592622305e+01 ppscbe1=-2.707617044e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.953629437e-01 lkt1=-7.824278632e-08 wkt1=-5.817825285e-08 pkt1=1.899607487e-13 kt2=-4.019094801e-02 lkt2=-5.623986592e-09 wkt2=-7.425247400e-09 pkt2=2.298378271e-14 at=1.619829214e+05 lat=-8.740708497e-02 wat=7.745375618e-03 pat=-3.079666683e-8 ute=-1.522233160e+00 lute=-6.183638592e-07 wute=-1.229961432e-06 pute=3.888438961e-12 ua1=1.248403606e-09 lua1=-1.804411272e-15 wua1=-3.603968216e-15 pua1=8.359019832e-21 ub1=-1.501811367e-18 lub1=1.884257516e-24 wub1=3.569488326e-24 pub1=-6.232784567e-30 uc1=3.168071888e-12 luc1=3.409463800e-17 wuc1=1.915102945e-17 puc1=1.049708130e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.22 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.233547157e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.274532987e-08 wvth0=-8.821092714e-08 pvth0=1.940783545e-13 k1=4.322980265e-01 lk1=2.290354845e-07 wk1=5.852102679e-07 pk1=-1.034063955e-12 k2=4.167122191e-03 lk2=-7.595777611e-08 wk2=-1.882744749e-07 pk2=3.376489246e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.489410334e+00 ldsub=2.580770446e-06 wdsub=6.924354866e-06 pdsub=-9.340265647e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.507121201e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.248992790e-08 wvoff=4.792095379e-08 pvoff=-1.208336804e-13 nfactor=2.535915471e+00 lnfactor=4.078665306e-07 wnfactor=2.176960983e-06 pnfactor=-3.863886733e-12 eta0=-2.287746183e-01 leta0=2.208577195e-07 weta0=1.136378997e-06 peta0=-1.094691106e-12 etab=8.131145842e-02 letab=4.133946247e-08 wetab=-4.058369249e-07 petab=-2.041860044e-13 u0=3.381781693e-02 lu0=-6.680492730e-09 wu0=-7.739682665e-10 pu0=-4.409137331e-15 ua=-3.458116995e-10 lua=-9.588258568e-16 wua=6.502986599e-16 pua=-1.075119411e-21 ub=1.130976655e-18 lub=1.021416273e-24 wub=-6.856039699e-25 pub=8.794109197e-31 uc=1.502659292e-10 luc=-1.324205014e-16 wuc=-2.857632557e-16 puc=4.528551467e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=6.427304155e+04 lvsat=3.107860877e-02 wvsat=5.923383665e-02 pvsat=-1.170541170e-7 a0=-6.103081915e-01 la0=2.601542635e-06 wa0=8.041458131e-06 pa0=-1.104799802e-11 ags=-4.217974222e-01 lags=1.756740021e-06 wags=1.688826944e-06 pags=-2.245630170e-12 a1=0.0 a2=0.42385546 b0=-6.155439406e-24 lb0=6.008546000e-30 wb0=3.050809353e-29 pb0=-2.978004839e-35 b1=0.0 keta=9.343023049e-02 lketa=-1.789801438e-07 wketa=-1.258512634e-07 pketa=2.342675965e-13 dwg=0.0 dwb=0.0 pclm=1.227253434e+00 lpclm=-1.672222791e-06 wpclm=-3.249432765e-06 ppclm=7.139976106e-12 pdiblc1=2.243127512e-01 lpdiblc1=3.274205370e-07 wpdiblc1=-1.755452639e-07 ppdiblc1=3.469013155e-13 pdiblc2=3.212200966e-03 lpdiblc2=4.346626400e-09 wpdiblc2=9.366012297e-09 ppdiblc2=-2.179673150e-14 pdiblcb=-4.944563519e-02 lpdiblcb=4.830789974e-08 wpdiblcb=6.779777293e-10 ppdiblcb=-1.339776198e-15 drout=8.528408000e-01 ldrout=-5.786932471e-7 pscbe1=5.784538022e+08 lpscbe1=4.621626191e+02 wpscbe1=1.703665918e+03 ppscbe1=-3.487396714e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-9.144845511e-06 lalpha0=1.813074251e-11 walpha0=2.704032152e-11 palpha0=-5.343535280e-17 alpha1=1.086627438e+00 lalpha1=-4.676079994e-07 walpha1=-1.337284493e-06 palpha1=2.642656028e-12 beta0=7.449738725e+00 lbeta0=1.266754807e-05 wbeta0=1.701998445e-05 pbeta0=-3.363380400e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.679801847e-01 lkt1=6.525875782e-08 wkt1=-5.825906639e-08 pkt1=1.901204472e-13 kt2=-7.282323658e-02 lkt2=5.886185362e-08 wkt2=7.557408473e-08 pkt2=-1.410341855e-13 at=1.771510203e+05 lat=-1.173813113e-01 wat=-4.068308861e-02 pat=6.490456476e-8 ute=-3.275796075e+00 lute=2.846914947e-06 wute=3.807485547e-06 pute=-6.066241361e-12 ua1=-2.531529433e-09 lua1=5.665250484e-15 wua1=5.963864993e-15 pua1=-1.054831981e-20 ub1=5.443922638e-19 lub1=-2.159319143e-24 wub1=1.901090271e-25 pub1=4.453285231e-31 uc1=-1.039974794e-10 luc1=2.458683418e-16 wuc1=6.134067940e-16 puc1=-1.069359396e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.23 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.841667251e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.099813825e-08 wvth0=2.621288451e-07 pvth0=-1.479009094e-13 k1=9.874452943e-01 lk1=-3.128637488e-07 wk1=-1.620513872e-06 pk1=1.119022784e-12 k2=-1.851773823e-01 lk2=1.088682111e-07 wk2=5.454289133e-07 pk2=-3.785453660e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.876654397e+00 ldsub=-7.049665158e-07 wdsub=-4.975986760e-06 pdsub=2.276086227e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-7.758134817e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.980105363e-08 wvoff=-1.502043658e-07 pvoff=7.256357659e-14 nfactor=3.264479119e+00 lnfactor=-3.033106744e-07 wnfactor=-3.970746006e-06 pnfactor=2.137111376e-12 eta0=-4.715281226e-01 leta0=4.578181542e-07 weta0=2.913868551e-08 peta0=-1.387397716e-14 etab=2.412787209e-01 letab=-1.148103413e-07 wetab=-1.198495941e-06 petab=5.695569972e-13 u0=2.766326795e-02 lu0=-6.728159131e-10 wu0=-1.219950617e-10 pu0=-5.045551847e-15 ua=-1.172891700e-09 lua=-1.514832936e-16 wua=-5.881447193e-16 pua=1.337697550e-22 ub=2.093119325e-18 lub=8.223417673e-26 wub=6.059720805e-25 pub=-3.813429598e-31 uc=-5.719003815e-11 luc=7.008473667e-17 wuc=3.877976020e-16 puc=-2.046318547e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.902380491e+04 lvsat=1.667985763e-02 wvsat=-1.531642220e-01 pvsat=9.027527433e-8 a0=2.583189677e+00 la0=-5.157455999e-07 wa0=-6.396882493e-06 pa0=3.045786043e-12 ags=1.407338691e+00 lags=-2.874558805e-08 wags=-7.365573499e-07 pags=1.218747529e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.738030033e-01 lketa=8.187583615e-08 wketa=3.177783144e-07 pketa=-1.987752051e-13 dwg=0.0 dwb=0.0 pclm=-1.385751826e+00 lpclm=8.784257117e-07 wpclm=8.102702856e-06 ppclm=-3.941252151e-12 pdiblc1=-2.765528811e-01 lpdiblc1=8.163335119e-07 wpdiblc1=2.991574971e-06 ppdiblc1=-2.744638762e-12 pdiblc2=9.419806541e-03 lpdiblc2=-1.712840875e-09 wpdiblc2=-1.199593703e-08 ppdiblc2=-9.445637253e-16 pdiblcb=2.389127038e-02 lpdiblcb=-2.327889391e-08 wpdiblcb=-1.355955459e-09 ppdiblcb=6.456192082e-16 drout=-2.494552533e-01 ldrout=4.972976131e-07 wdrout=-5.771431887e-07 pdrout=5.633702437e-13 pscbe1=1.291806799e+09 lpscbe1=-2.341669223e+02 wpscbe1=-3.648774159e+03 ppscbe1=1.737312733e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.289806226e-05 lalpha0=-1.314749331e-11 walpha0=-7.647496508e-11 palpha0=4.760964499e-17 alpha1=3.767451235e-01 lalpha1=2.253336839e-07 walpha1=2.674568986e-06 palpha1=-1.273458578e-12 beta0=3.253329128e+01 lbeta0=-1.181741058e-05 wbeta0=-6.304794120e-05 pbeta0=4.452338067e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.236107223e-01 lkt1=2.194812831e-08 wkt1=2.712027395e-07 pkt1=-1.314790822e-13 kt2=9.325787446e-03 lkt2=-2.132676610e-08 wkt2=-1.304250988e-07 pkt2=6.004903355e-14 at=4.960931399e+04 lat=7.116739710e-03 wat=1.009528817e-01 pat=-7.335140480e-8 ute=1.007947713e+00 lute=-1.334601580e-06 wute=-6.225017667e-06 pute=3.726846196e-12 ua1=5.416821995e-09 lua1=-2.093421486e-15 wua1=-9.514190675e-15 pua1=4.560367534e-21 ub1=-1.388221491e-18 lub1=-2.728252830e-25 wub1=-2.629157462e-24 pub1=3.197316037e-30 uc1=3.920554572e-10 luc1=-2.383467875e-16 wuc1=-1.393195215e-15 puc1=8.893570623e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.24 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.462432295e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.617232026e-08 wvth0=-9.127629017e-08 pvth0=2.036799811e-14 k1=-4.462581406e-02 lk1=1.785424604e-07 wk1=1.298853683e-06 pk1=-2.709932064e-13 k2=1.575393653e-01 lk2=-5.431157018e-08 wk2=-4.530767430e-07 pk2=9.687912315e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.153734590e-01 ldsub=3.841554494e-08 wdsub=-6.085653180e-07 pdsub=1.965996510e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.400137708e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.472967018e-11 wvoff=1.676737799e-08 pvoff=-6.937681634e-15 nfactor=2.495136391e+00 lnfactor=6.300109494e-08 wnfactor=3.109409937e-07 pnfactor=9.844605514e-14 eta0=0.49 etab=1.910278903e-03 letab=-8.384087608e-10 wetab=-7.494999385e-09 petab=2.478572728e-15 u0=3.357104954e-02 lu0=-3.485723408e-09 wu0=-1.613181330e-08 pu0=2.577298969e-15 ua=-8.915624399e-10 lua=-2.854342821e-16 wua=-7.509814663e-16 pua=2.113021923e-22 ub=1.924065949e-18 lub=1.627265745e-25 wub=1.618320143e-25 pub=-1.698718852e-31 uc=1.640827545e-10 luc=-3.527120574e-17 wuc=-2.572489332e-16 puc=1.024980224e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.165365894e+05 lvsat=-1.181329507e-03 wvsat=-3.530647615e-02 pvsat=3.415895867e-8 a0=1.5 ags=2.547688899e+00 lags=-5.717073745e-07 wags=-9.153052131e-07 pags=2.069830455e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.560495070e-02 lketa=-8.308109442e-09 wketa=-1.396456155e-07 pketa=1.902079523e-14 dwg=0.0 dwb=0.0 pclm=3.506056264e-01 lpclm=5.168341970e-08 wpclm=3.563941332e-07 ppclm=-2.529557012e-13 pdiblc1=1.826620147e+00 lpdiblc1=-1.850628808e-07 wpdiblc1=-3.000380505e-06 ppdiblc1=1.083469502e-13 pdiblc2=8.864730888e-03 lpdiblc2=-1.448549374e-09 wpdiblc2=-2.695224928e-08 ppdiblc2=6.176674961e-15 pdiblcb=-2.924087145e-01 lpdiblcb=1.273229157e-07 wpdiblcb=1.325352999e-06 ppdiblcb=-6.310482753e-13 drout=6.095479465e-01 ldrout=8.829526556e-08 wdrout=1.154286377e-06 pdrout=-2.610257043e-13 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.465450645e-05 lalpha0=4.732636541e-12 walpha0=5.274076208e-11 palpha0=-1.391461447e-17 alpha1=0.85 beta0=-3.230690459e+00 lbeta0=5.211108629e-06 wbeta0=5.985155848e-05 pbeta0=-1.399349550e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.446665968e-01 lkt1=-1.564001184e-08 wkt1=-1.899183510e-07 pkt1=8.807726938e-14 kt2=-3.116452394e-02 lkt2=-2.047871194e-09 wkt2=-7.000030631e-08 pkt2=3.127861454e-14 at=9.235246539e+04 lat=-1.323481343e-02 wat=-7.136271010e-02 pat=8.694251837e-9 ute=-2.354879333e+00 lute=2.665614384e-07 wute=6.567354300e-07 pute=4.501958030e-13 ua1=1.356030169e-09 lua1=-1.599323086e-16 wua1=-4.530399546e-15 pua1=2.187405161e-21 ub1=-3.727401675e-18 lub1=8.409426132e-25 wub1=1.162068866e-23 pub1=-3.587548696e-30 uc1=-3.170077008e-10 luc1=9.926370828e-17 wuc1=1.094375105e-15 puc1=-2.950647196e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.25 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='7.832310539e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.715019890e-08 wvth0=-4.870291161e-07 pvth0=1.098619591e-13 k1=4.931050082e-01 lk1=5.694216317e-08 wk1=-2.708135376e-10 pk1=2.278561067e-14 k2=-3.118944394e-02 lk2=-1.163319218e-08 wk2=8.499234707e-08 pk2=-2.479766861e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.949779736e-01 ldsub=-9.265390157e-08 wdsub=-1.931363806e-07 pdsub=1.026562128e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-5.638404937e-03 lcdscd=2.496180739e-09 wcdscd=5.470944770e-08 pcdscd=-1.237177566e-14 cit=0.0 voff='-2.446740146e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.359271923e-08 wvoff=5.384288674e-07 pvoff=-1.249041242e-13 nfactor=-1.540586399e+00 lnfactor=9.756233037e-07 wnfactor=1.747296423e-05 pnfactor=-3.782505231e-12 eta0=1.377471867e+00 leta0=-2.006893380e-07 weta0=6.028800406e-07 peta0=-1.363328809e-13 etab=-3.521303131e-02 letab=7.556508117e-09 wetab=4.354878357e-07 petab=-9.769579367e-14 u0=-4.339233702e-03 lu0=5.087156403e-09 wu0=-1.524974200e-08 pu0=2.377830894e-15 ua=-6.749666627e-09 lua=1.039293966e-15 wua=7.792177348e-15 pua=-1.720613569e-21 ub=7.661363531e-18 lub=-1.134682951e-24 wub=-1.347426977e-23 pub=2.913741628e-30 uc=-2.264736401e-10 luc=5.304765511e-17 wuc=9.862569928e-16 puc=-1.787034337e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.109476091e+05 lvsat=8.254013386e-05 wvsat=1.084669381e-01 pvsat=1.646613870e-9 a0=1.5 ags=-2.725045681e+00 lags=6.206477325e-07 wags=-5.916754457e-12 pags=9.238183736e-19 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=7.781446191e-03 lketa=-6.538933426e-09 wketa=-6.967213643e-08 pketa=3.197272573e-15 dwg=0.0 dwb=0.0 pclm=5.388206768e-01 lpclm=9.121221069e-09 wpclm=-2.077578437e-07 ppclm=-1.253806297e-13 pdiblc1=2.359042693e+00 lpdiblc1=-3.054627857e-07 wpdiblc1=-7.843734467e-06 ppdiblc1=1.203603642e-12 pdiblc2=-1.570608770e-02 lpdiblc2=4.107797258e-09 wpdiblc2=1.565499552e-08 ppdiblc2=-3.458356948e-15 pdiblcb=1.120676856e+00 lpdiblcb=-1.922266030e-07 wpdiblcb=-4.780721519e-06 ppdiblcb=7.497549918e-13 drout=4.516027116e-01 ldrout=1.240123692e-07 wdrout=4.896295556e-06 pdrout=-1.107228692e-12 pscbe1=7.850767286e+08 lpscbe1=3.374688911e+00 wpscbe1=1.006949609e+02 ppscbe1=-2.277075567e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.083252961e-05 lalpha0=-1.030899845e-12 walpha0=-7.058061165e-13 palpha0=-1.828421326e-18 alpha1=1.837382488e+00 lalpha1=-2.232827263e-07 walpha1=-2.918981076e-06 palpha1=6.600867046e-13 beta0=9.327764020e+00 lbeta0=2.371189967e-06 wbeta0=6.112838551e-05 pbeta0=-1.428223206e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.331906060e-01 lkt1=4.378453513e-09 wkt1=2.874000947e-07 pkt1=-1.986161466e-14 kt2=-2.650655854e-02 lkt2=-3.101204857e-09 wkt2=1.053719629e-07 pkt2=-8.379368922e-15 at=1.150888746e+05 lat=-1.837633407e-02 wat=-6.228187239e-01 pat=1.333983090e-7 ute=1.987849026e+00 lute=-7.154857818e-07 wute=1.418809837e-07 pute=5.666229281e-13 ua1=5.008738400e-09 lua1=-9.859411372e-16 wua1=8.159284493e-15 pua1=-6.821892292e-22 ub1=-2.016597456e-18 lub1=4.540681903e-25 wub1=-1.249786236e-23 pub1=1.866523956e-30 uc1=3.321514218e-10 luc1=-4.753453906e-17 wuc1=-1.467657294e-15 puc1=2.843030389e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.26 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.304860242e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.768760094e-08 wvth0=5.131328281e-07 pvth0=-4.629932617e-14 k1=7.069074261e-01 lk1=2.355990885e-08 wk1=5.917473316e-07 pk1=-6.964973445e-14 k2=-1.005113253e-01 lk2=-8.095509190e-10 wk2=-9.690911799e-08 pk2=3.603698539e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.289742177e-01 ldsub=-4.280339138e-09 wdsub=3.833604585e-07 pdsub=1.264430231e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=3.060418107e-02 lcdscd=-3.162591669e-09 wcdscd=-8.440829895e-08 pcdscd=9.349512825e-15 cit=0.0 voff='9.710513754e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.977131047e-08 wvoff=-8.252317455e-07 pvoff=8.801238925e-14 nfactor=9.877720445e+00 lnfactor=-8.071854536e-07 wnfactor=-3.245888202e-05 pnfactor=4.013653515e-12 eta0=4.763329940e-01 leta0=-5.998911901e-08 weta0=-1.406122568e-06 peta0=1.773447504e-13 etab=1.500326779e-01 letab=-2.136701594e-08 wetab=-5.947852485e-07 petab=6.316692461e-14 u0=1.635267749e-01 lu0=-2.112277071e-08 wu0=-3.762372093e-07 pu0=5.874097009e-14 ua=1.697280683e-08 lua=-2.664638150e-15 wua=-5.375949692e-14 pua=7.889818645e-21 ub=-1.396242758e-17 lub=2.241569298e-24 wub=5.054657819e-23 pub=-7.082217490e-30 uc=5.266491414e-10 luc=-6.454192351e-17 wuc=-1.380318047e-15 puc=1.908041267e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-9.405219098e+04 lvsat=3.209038892e-02 wvsat=5.492619481e-01 pvsat=-6.717735582e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.519339594e-01 lketa=-9.150073022e-08 wketa=-2.641277947e-06 pketa=4.047175174e-13 dwg=0.0 dwb=0.0 pclm=2.605040018e+00 lpclm=-3.134900019e-07 wpclm=-5.756253401e-06 ppclm=7.409392726e-13 pdiblc1=7.311991496e-01 lpdiblc1=-5.129780627e-08 wpdiblc1=-1.106320543e-06 ppdiblc1=1.516507813e-13 pdiblc2=1.462683294e-02 lpdiblc2=-6.282636394e-10 wpdiblc2=-1.839020505e-08 ppdiblc2=1.857324488e-15 pdiblcb=-8.436781848e-01 lpdiblcb=1.144799357e-07 wpdiblcb=2.188779206e-06 ppdiblcb=-3.384349734e-13 drout=4.635200135e+00 ldrout=-5.291977980e-07 wdrout=-1.221498318e-05 pdrout=1.564457925e-12 pscbe1=8.624336049e+08 lpscbe1=-8.703504333e+00 wpscbe1=-2.099365967e+02 ppscbe1=2.573001320e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.188879730e-05 lalpha0=-2.757181256e-12 walpha0=-6.462076899e-11 palpha0=8.151005317e-18 alpha1=-1.453892472e+00 lalpha1=2.906037808e-07 walpha1=6.810955844e-06 palpha1=-8.591067263e-13 beta0=6.931149233e+01 lbeta0=-6.994429437e-06 wbeta0=-1.579296821e-04 pbeta0=1.992061838e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-6.425863786e-01 lkt1=5.268627187e-08 wkt1=1.157755826e-06 pkt1=-1.557554772e-13 kt2=-1.167450682e-01 lkt2=1.098827508e-08 wkt2=2.597570561e-07 pkt2=-3.248443984e-14 at=-2.489356391e+05 lat=3.846099742e-02 wat=1.146221855e+00 pat=-1.428126109e-7 ute=-2.170141203e+01 lute=2.983260683e-06 wute=6.025603010e-05 pute=-8.819359858e-12 ua1=-2.584295612e-08 lua1=3.831119038e-15 wua1=7.632856654e-14 pua1=-1.132586825e-20 ub1=1.540697490e-17 lub1=-2.266378703e-24 wub1=-4.345504462e-23 pub1=6.700054566e-30 uc1=-4.011452666e-10 luc1=6.695947268e-17 wuc1=1.621022593e-15 puc1=-1.979510838e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.27 nmos lmin=2.0e-05 lmax=0.0001 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.190746862e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.108125260e-08 wvth0=-2.129199822e-09 pvth0=4.253318521e-14 k1=5.344591002e-01 lk1=3.397603097e-07 wk1=1.111346905e-08 pk1=-2.220041692e-13 k2=-2.587186719e-02 lk2=-7.955865334e-08 wk2=-2.103903829e-10 pk2=4.202786903e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.080533089e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.604577012e-08 wvoff=8.586471678e-09 pvoff=-1.715245260e-13 nfactor=2.419326758e+00 lnfactor=5.891426789e-06 wnfactor=5.728458176e-07 pnfactor=-1.144324596e-11 eta0=0.08 etab=-0.07 u0=3.331007502e-02 lu0=-4.923268569e-08 wu0=-3.532766031e-09 pu0=7.057101470e-14 ua=-8.605860935e-10 lua=3.112478025e-15 wua=2.615327364e-16 pua=-5.224413510e-21 ub=1.916544460e-18 lub=-7.475558700e-24 wub=-6.191158015e-25 pub=1.236754145e-29 uc=4.982766889e-11 luc=4.223820340e-16 wuc=-1.777224155e-17 puc=3.550207143e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.253958055e+00 la0=3.361822778e-06 wa0=1.737682905e-07 pa0=-3.471219004e-12 ags=4.144789130e-01 lags=1.272653665e-08 wags=-3.486438228e-08 pags=6.964556420e-13 a1=0.0 a2=0.42385546 b0=-5.261963924e-25 lb0=5.260708209e-29 b1=7.785514628e-24 lb1=-1.555244990e-28 wb1=-1.523066213e-29 pb1=3.042497780e-34 keta=-1.595293910e-02 lketa=2.056551011e-07 wketa=1.884659271e-08 pketa=-3.764820991e-13 dwg=0.0 dwb=0.0 pclm=-1.115928690e-01 lpclm=3.897820945e-06 wpclm=3.654620441e-07 ppclm=-7.300519495e-12 pdiblc1=0.39 pdiblc2=2.932071753e-03 lpdiblc2=-9.379484098e-09 wpdiblc2=8.689549233e-10 ppdiblc2=-1.735836173e-14 pdiblcb=5.959123923e-01 lpdiblcb=-6.207642177e-05 wpdiblcb=-1.942890293e-22 ppdiblcb=9.769962617e-27 drout=0.56 pscbe1=8.920131824e+08 lpscbe1=-1.967597506e+03 wpscbe1=-4.346853224e+02 ppscbe1=8.683333118e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.844064645e-01 lkt1=-6.379086479e-07 wkt1=-8.217583833e-08 pkt1=1.641555722e-12 kt2=-4.589540693e-02 lkt2=9.655954614e-08 wkt2=-1.417775330e-09 pkt2=2.832167281e-14 at=140000.0 ute=-1.647300853e+00 lute=-2.856570414e-06 wute=-5.080880770e-07 pute=1.014963653e-11 ua1=6.731339193e-10 lua1=-6.836910839e-15 wua1=-8.450306964e-16 pua1=1.688044812e-20 ub1=-1.039765919e-18 lub1=1.227745143e-23 wub1=1.024632243e-24 pub1=-2.046819303e-29 uc1=1.306819906e-11 luc1=4.193256512e-17 wuc1=8.652776088e-18 puc1=-1.728490319e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.28 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.5216318+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.029854552 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.71425 eta0=0.08 etab=-0.07 u0=0.0308455 ua=-7.0477628e-10 ub=1.54232e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.42225 ags=0.415116 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.29 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.137418539e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.293128287e-8 k1=5.483309743e-01 lk1=2.501663785e-8 k2=-2.596763155e-02 lk2=-3.100260617e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077791411e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.619850412e-8 nfactor=2.647232228e+00 lnfactor=5.345428661e-7 eta0=0.08 etab=-0.07 u0=3.099400868e-02 lu0=-1.184525426e-9 ua=-7.496494897e-10 lua=3.579148231e-16 ub=1.611793036e-18 lub=-5.541263855e-25 uc=8.123639508e-11 luc=-8.187021115e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.561973407e+00 la0=-1.114452897e-6 ags=4.088306236e-01 lags=5.013301686e-8 a1=0.0 a2=0.42385546 b0=4.202027848e-24 lb0=-1.670783420e-29 b1=0.0 keta=-1.059979967e-02 lketa=3.941726389e-8 dwg=0.0 dwb=0.0 pclm=-3.193698668e-01 lpclm=3.213592108e-06 wpclm=1.110223025e-22 ppclm=-1.332267630e-27 pdiblc1=0.39 pdiblc2=1.440006234e-03 lpdiblc2=8.155846848e-9 pdiblcb=-4.983398045e+00 lpdiblcb=1.971526497e-5 drout=0.56 pscbe1=7.870702449e+08 lpscbe1=5.141046490e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141332445e-01 lkt1=-1.760138183e-8 kt2=-3.996812420e-02 lkt2=-8.722206193e-9 at=140000.0 ute=-1.817437128e+00 lute=2.164494252e-7 ua1=3.748619787e-10 lua1=-3.508062434e-16 ub1=-4.991379884e-19 lub1=5.900584965e-25 uc1=3.254985601e-12 luc1=9.501449495e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.30 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.259943688e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.421361748e-8 k1=5.402698164e-01 lk1=5.706889798e-8 k2=-2.744592236e-02 lk2=-2.512472084e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064515944e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.091999792e-8 nfactor=2.746465137e+00 lnfactor=1.399793225e-7 eta0=0.08 etab=-0.07 u0=3.195628193e-02 lu0=-5.010654727e-9 ua=-5.258090296e-10 lua=-5.321052884e-16 ub=1.379512085e-18 lub=3.694542658e-25 uc=5.722333245e-11 luc=1.360899167e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.031231535e+00 la0=9.958489658e-7 ags=1.915997610e-01 lags=9.138724701e-7 a1=0.0 a2=0.42385546 b0=-2.082155696e-24 lb0=8.278934222e-30 b1=0.0 keta=-1.749000880e-03 lketa=4.225284179e-09 pketa=-1.734723476e-30 dwg=0.0 dwb=0.0 pclm=4.738214857e-01 lpclm=5.975541666e-8 pdiblc1=0.39 pdiblc2=2.149708243e-03 lpdiblc2=5.333975140e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.082391335e+08 lpscbe1=-3.275991519e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.150424779e-01 lkt1=-1.398614617e-8 kt2=-4.270263241e-02 lkt2=2.150570337e-9 at=1.646028932e+05 lat=-9.782444936e-2 ute=-1.938283263e+00 lute=6.969500930e-7 ua1=2.931550244e-11 lua1=1.023133540e-15 ub1=-2.943865257e-19 lub1=-2.240611654e-25 uc1=9.646151264e-12 luc1=6.960235108e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.31 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.935162473e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.839480260e-8 k1=6.302528454e-01 lk1=-1.207498050e-7 k2=-5.951911442e-02 lk2=3.825626861e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.886133968e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.336345769e-8 nfactor=3.272300222e+00 lnfactor=-8.991423180e-7 eta0=1.556200357e-01 leta0=-1.494354750e-7 etab=-5.596804500e-02 letab=-2.772905143e-8 u0=3.355601231e-02 lu0=-8.171939531e-9 ua=-1.258399038e-10 lua=-1.322498677e-15 ub=8.990623895e-19 lub=1.318888206e-24 uc=5.360287210e-11 luc=2.076351371e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.430964044e+04 lvsat=-8.516435621e-3 a0=2.109817335e+00 la0=-1.135583262e-6 ags=1.494697789e-01 lags=9.971270444e-7 a1=0.0 a2=0.42385546 b0=4.164311393e-24 lb0=-4.064934266e-30 b1=0.0 keta=5.085943942e-02 lketa=-9.973614859e-08 wketa=-1.994931997e-23 pketa=-4.423544864e-29 dwg=0.0 dwb=0.0 pclm=1.280914582e-01 lpclm=7.429649702e-7 pdiblc1=1.649323322e-01 lpdiblc1=4.447643207e-7 pdiblc2=6.380373791e-03 lpdiblc2=-3.026395354e-9 pdiblcb=-4.921630060e-02 lpdiblcb=4.785470340e-8 drout=8.528408000e-01 ldrout=-5.786932471e-7 pscbe1=1.154740475e+09 lpscbe1=-7.174936905e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.887283200e-09 lalpha0=5.555455173e-14 alpha1=6.342739440e-01 lalpha1=4.263040254e-7 beta0=1.320696502e+01 lbeta0=1.290485941e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.876870551e-01 lkt1=1.295694180e-7 kt2=-4.725934087e-02 lkt2=1.115524596e-8 at=1.633894479e+05 lat=-9.542651645e-2 ute=-1.987865646e+00 lute=7.949316238e-7 ua1=-5.141762198e-10 lua1=2.097147098e-15 pua1=8.271806126e-37 ub1=6.086990610e-19 lub1=-2.008681104e-24 pub1=-7.703719778e-46 uc1=1.034951732e-10 luc1=-1.158560798e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.32 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.728351421e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.687738636e-10 k1=4.392858589e-01 lk1=6.565994532e-8 k2=-6.791127560e-04 lk2=-1.917957525e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.934635650e-01 ldsub=6.494860950e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.283898860e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.255500608e-9 nfactor=1.921323762e+00 lnfactor=4.195944397e-7 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=1.977584763e-22 peta0=-7.285838599e-29 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.762200157e-02 lu0=-2.379538021e-9 ua=-1.371839134e-09 lua=-1.062339720e-16 ub=2.298097091e-18 lub=-4.675993133e-26 uc=7.398743477e-11 luc=8.654082393e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.721405808e+04 lvsat=4.721661776e-2 a0=4.193627844e-01 la0=5.145302813e-7 ags=1.158188796e+00 lags=1.248009777e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.631044528e-02 lketa=1.463759397e-8 dwg=0.0 dwb=0.0 pclm=1.355090508e+00 lpclm=-4.547529740e-7 pdiblc1=7.353854155e-01 lpdiblc1=-1.120754702e-7 pdiblc2=5.362028211e-03 lpdiblc2=-2.032351573e-9 pdiblcb=2.343260119e-02 lpdiblcb=-2.306050500e-08 wpdiblcb=3.903127821e-24 ppdiblcb=-2.385244779e-30 drout=-4.446812800e-01 ldrout=6.878647659e-07 pdrout=2.220446049e-28 pscbe1=5.756251585e+07 lpscbe1=3.535012140e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.970567686e-06 lalpha0=2.957074856e-12 walpha0=-5.293955920e-28 palpha0=-6.882142696e-34 alpha1=1.281452112e+00 lalpha1=-2.054298828e-7 beta0=1.120652299e+01 lbeta0=3.243189417e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.318729451e-01 lkt1=-2.252634408e-8 kt2=-3.479216166e-02 lkt2=-1.014416479e-9 at=8.375791069e+04 lat=-1.769530623e-2 ute=-1.097743715e+00 lute=-7.394843689e-8 ua1=2.198525948e-09 lua1=-5.508191447e-16 ub1=-2.277567454e-18 lub1=8.087075466e-25 uc1=-7.921055025e-11 luc1=6.248955431e-17 puc1=-1.292469707e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.33 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.153678631e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.928258575e-8 k1=3.947279698e-01 lk1=8.687556041e-8 k2=4.280392337e-03 lk2=-2.154097416e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.095184973e-01 ldsub=1.049178783e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.343419918e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.421488753e-9 nfactor=2.600316138e+00 lnfactor=9.630172565e-8 eta0=0.49 etab=-0.000625 u0=2.811425844e-02 lu0=-2.613919240e-09 wu0=2.775557562e-23 ua=-1.145591476e-09 lua=-2.139586271e-16 ub=1.978807687e-18 lub=1.052652480e-25 uc=7.706502979e-11 luc=-5.999455450e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.045937246e+05 lvsat=1.037337287e-2 a0=1.5 ags=2.238075265e+00 lags=-5.016927259e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.163195547e-02 lketa=-1.874083449e-9 dwg=0.0 dwb=0.0 pclm=4.711604765e-01 lpclm=-3.388206463e-8 pdiblc1=8.117032664e-01 lpdiblc1=-1.484131464e-7 pdiblc2=-2.522103509e-04 lpdiblc2=6.407895190e-10 pdiblcb=1.559088000e-01 lpdiblcb=-8.613719240e-08 ppdiblcb=2.081668171e-29 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.185727360e-06 lalpha0=2.584115772e-14 alpha1=0.85 beta0=1.701486070e+01 lbeta0=4.776307318e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.089088954e-01 lkt1=1.415324515e-8 kt2=-5.484301818e-02 lkt2=8.532518139e-9 at=6.821312074e+04 lat=-1.029387212e-2 ute=-2.132730218e+00 lute=4.188458967e-7 ua1=-1.764351194e-10 lua1=5.799853180e-16 ub1=2.034441167e-19 lub1=-3.725913786e-25 pub1=1.925929944e-46 uc1=5.317860243e-11 luc1=-5.456872969e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.34 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.974970253e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.372254007e-09 wvth0=3.576812492e-07 pvth0=-8.088460698e-14 k1=4.930134021e-01 lk1=6.464968589e-8 k2=-5.131989890e-03 lk2=-1.941249570e-08 wk2=7.959164690e-09 pk2=-1.799853666e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.296255798e-01 ldsub=-5.792425694e-08 wdsub=6.372491664e-11 pdsub=-1.441049775e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.286776183e-02 lcdscd=-1.688729789e-09 wcdscd=1.387778781e-23 cit=0.0 voff='-1.737695956e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.494511867e-09 wvoff=3.288154100e-07 pvoff=-7.435700155e-14 nfactor=5.138848303e+00 lnfactor=-4.777517840e-07 wnfactor=-2.273328352e-06 pnfactor=5.140813803e-13 eta0=1.581403705e+00 leta0=-2.468056683e-07 weta0=1.573773112e-14 peta0=-3.558867867e-21 etab=1.433521275e-01 letab=-3.255841171e-08 wetab=-9.240112913e-08 petab=2.089522174e-14 u0=-8.717456487e-03 lu0=5.715057447e-09 wu0=-2.306480789e-09 pu0=5.215783396e-16 ua=-4.117754007e-09 lua=4.581543190e-16 wua=1.150144447e-17 pua=-2.600890647e-24 ub=2.543297387e-18 lub=-2.238619480e-26 wub=1.656177044e-24 pub=-3.745212521e-31 uc=2.061964889e-10 luc=-2.980121719e-17 wuc=-2.928379216e-16 puc=6.622119624e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.280291486e+05 lvsat=-1.753982017e-02 wvsat=-2.376591097e-01 pvsat=5.374328043e-8 a0=1.5 ags=-2.725047683e+00 lags=6.206480450e-07 wags=-3.330669074e-22 pags=4.163336342e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.859815628e-01 lketa=-7.369793403e-08 wketa=-8.921101337e-07 pketa=2.017382172e-13 dwg=0.0 dwb=0.0 pclm=2.289816123e-02 lpclm=6.748618229e-08 wpclm=1.317454603e-06 ppclm=-2.979239140e-13 pdiblc1=-2.942002886e-01 lpdiblc1=1.016714599e-07 ppdiblc1=5.551115123e-29 pdiblc2=-1.041058628e-02 lpdiblc2=2.937964019e-09 ppdiblc2=-8.673617380e-31 pdiblcb=-4.964630236e-01 lpdiblcb=6.138756232e-8 drout=2.107836980e+00 ldrout=-2.505218234e-7 pscbe1=8.191380802e+08 lpscbe1=-4.327808912e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.059378171e-05 lalpha0=-1.649386622e-12 alpha1=0.85 beta0=2.830344734e+01 lbeta0=-2.075125096e-06 wbeta0=5.030914472e-06 pbeta0=-1.137670875e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.923387179e-01 lkt1=-1.220746851e-08 wkt1=-1.289978070e-07 pkt1=2.917104808e-14 kt2=9.136848570e-03 lkt2=-5.935633008e-9 at=-1.610402072e+05 lat=4.154855845e-02 wat=1.934967105e-01 pat=-4.375657212e-8 ute=2.035842074e+00 lute=-5.238183671e-7 ua1=7.768720193e-09 lua1=-1.216700324e-15 ub1=-6.244158411e-18 lub1=1.085443667e-24 uc1=-1.643023312e-10 luc1=4.863458112e-17 puc1=-2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.35 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=2.0e-06 wmax=3.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='1.176143311e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-9.858886246e-08 wvth0=-1.395612187e-06 pvth0=1.928676170e-13 k1=0.90707349 k2=-1.372151317e-01 lk2=1.210437729e-09 wk2=1.159768416e-08 pk2=-2.367957542e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587010672e-01 ldsub=-9.587241274e-12 wdsub=-1.486914722e-10 pdsub=1.875534753e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.321743718e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-1.474168590e-7 nfactor=-8.343868507e+00 lnfactor=1.627385688e-06 wnfactor=2.140927341e-05 pnfactor=-3.183625328e-12 eta0=6.941575510e-04 leta0=-2.367699262e-15 weta0=-3.672137572e-14 peta0=4.631887448e-21 etab=-6.517384797e-02 wetab=4.142593021e-8 u0=5.160786376e-02 lu0=-3.703896755e-09 wu0=-4.537334693e-08 pu0=7.245866552e-15 ua=-1.262823224e-09 lua=1.239684637e-17 wua=1.501679709e-16 pua=-2.425172742e-23 ub=5.317291396e-18 lub=-4.555065233e-25 wub=-6.449707982e-24 pub=8.910992123e-31 uc=1.532944232e-11 wuc=1.312871760e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.165870995e+04 lvsat=2.769088331e-02 wvsat=4.534976832e-01 pvsat=-5.417117659e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.045636319e+00 lketa=1.342155556e-07 wketa=2.081590312e-06 pketa=-2.625634756e-13 dwg=0.0 dwb=0.0 pclm=1.645277110e+00 lpclm=-1.858255773e-07 wpclm=-2.918923594e-06 ppclm=3.635272321e-13 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.986056660e+01 lbeta0=-7.568874690e-07 wbeta0=-1.173880043e-05 pbeta0=1.480685332e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705235600e-01 wkt1=5.783321264e-8 kt2=-0.028878939 at=2.915115102e+05 lat=-2.911105650e-02 wat=-4.514923244e-01 pat=5.694943583e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.36 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.179862952e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.282310025e-08 wvth0=8.881784197e-22 k1=5.401400138e-01 lk1=2.262776067e-7 k2=-2.597941323e-02 lk2=-7.741029901e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.036641300e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.163306452e-8 nfactor=2.712150501e+00 lnfactor=4.193987468e-8 eta0=0.08 etab=-0.07 u0=3.150421777e-02 lu0=-1.315863568e-8 ua=-7.268974247e-10 lua=4.418949960e-16 ub=1.600068716e-18 lub=-1.153596196e-24 uc=4.074296558e-11 luc=6.038593027e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.342783843e+00 la0=1.587426753e-6 ags=3.966571561e-01 lags=3.687363767e-7 a1=0.0 a2=0.42385546 b0=-5.261963924e-25 lb0=5.260708209e-29 b1=0.0 keta=-6.319055684e-03 lketa=1.320733586e-8 dwg=0.0 dwb=0.0 pclm=7.522173340e-02 lpclm=1.659870397e-7 pdiblc1=0.39 pdiblc2=3.376258697e-03 lpdiblc2=-1.825262290e-8 pdiblcb=5.959123923e-01 lpdiblcb=-6.207642177e-05 wpdiblcb=-1.665334537e-22 ppdiblcb=2.930988785e-26 drout=0.56 pscbe1=6.698134574e+08 lpscbe1=2.471094420e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.264125957e-01 lkt1=2.012115416e-7 kt2=-4.662013646e-02 lkt2=1.110368417e-7 at=140000.0 ute=-1.907022139e+00 lute=2.331657318e-6 ua1=2.411764120e-10 lua1=1.791931074e-15 ub1=-5.160008166e-19 lub1=1.814648506e-24 wub1=7.703719778e-40 uc1=1.749127103e-11 luc1=-4.642332218e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.37 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.5216318+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.55146741 k2=-0.029854552 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.71425 eta0=0.08 etab=-0.07 u0=0.0308455 ua=-7.0477628e-10 ub=1.54232e-18 uc=7.0972e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.42225 ags=0.415116 a1=0.0 a2=0.42385546 b0=2.1073e-24 b1=0.0 keta=-0.0056579 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0024625373 pdiblcb=-2.5116166 drout=0.56 pscbe1=793515780.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.31634 kt2=-0.041061662 at=140000.0 ute=-1.7903 ua1=3.3088e-10 ub1=-4.2516e-19 uc1=1.5167332e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.38 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.137418539e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.293128287e-8 k1=5.483309743e-01 lk1=2.501663785e-8 k2=-2.596763155e-02 lk2=-3.100260617e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.077791411e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.619850412e-8 nfactor=2.647232228e+00 lnfactor=5.345428661e-7 eta0=0.08 etab=-0.07 u0=3.099400868e-02 lu0=-1.184525426e-9 ua=-7.496494897e-10 lua=3.579148231e-16 ub=1.611793036e-18 lub=-5.541263855e-25 uc=8.123639508e-11 luc=-8.187021115e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.561973407e+00 la0=-1.114452897e-6 ags=4.088306236e-01 lags=5.013301686e-8 a1=0.0 a2=0.42385546 b0=4.202027848e-24 lb0=-1.670783420e-29 b1=0.0 keta=-1.059979967e-02 lketa=3.941726389e-8 dwg=0.0 dwb=0.0 pclm=-3.193698668e-01 lpclm=3.213592108e-06 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=1.440006234e-03 lpdiblc2=8.155846848e-9 pdiblcb=-4.983398045e+00 lpdiblcb=1.971526497e-5 drout=0.56 pscbe1=7.870702449e+08 lpscbe1=5.141046490e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.141332445e-01 lkt1=-1.760138183e-8 kt2=-3.996812420e-02 lkt2=-8.722206193e-9 at=140000.0 ute=-1.817437128e+00 lute=2.164494252e-7 ua1=3.748619787e-10 lua1=-3.508062434e-16 ub1=-4.991379884e-19 lub1=5.900584965e-25 uc1=3.254985601e-12 luc1=9.501449495e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.39 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.259943688e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.421361748e-8 k1=5.402698164e-01 lk1=5.706889798e-8 k2=-2.744592236e-02 lk2=-2.512472084e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.064515944e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.091999792e-8 nfactor=2.746465137e+00 lnfactor=1.399793225e-7 eta0=0.08 etab=-0.07 u0=3.195628193e-02 lu0=-5.010654727e-9 ua=-5.258090296e-10 lua=-5.321052884e-16 ub=1.379512085e-18 lub=3.694542658e-25 uc=5.722333245e-11 luc=1.360899167e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.031231535e+00 la0=9.958489658e-7 ags=1.915997610e-01 lags=9.138724701e-7 a1=0.0 a2=0.42385546 b0=-2.082155696e-24 lb0=8.278934222e-30 b1=0.0 keta=-1.749000880e-03 lketa=4.225284179e-09 wketa=1.734723476e-24 dwg=0.0 dwb=0.0 pclm=4.738214857e-01 lpclm=5.975541666e-8 pdiblc1=0.39 pdiblc2=2.149708243e-03 lpdiblc2=5.333975140e-9 pdiblcb=-0.025 drout=0.56 pscbe1=8.082391335e+08 lpscbe1=-3.275991519e+1 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.150424779e-01 lkt1=-1.398614617e-8 kt2=-4.270263241e-02 lkt2=2.150570337e-9 at=1.646028932e+05 lat=-9.782444936e-2 ute=-1.938283263e+00 lute=6.969500930e-7 ua1=2.931550244e-11 lua1=1.023133540e-15 ub1=-2.943865257e-19 lub1=-2.240611654e-25 uc1=9.646151264e-12 luc1=6.960235108e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.40 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.935162473e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.839480260e-8 k1=6.302528454e-01 lk1=-1.207498050e-7 k2=-5.951911442e-02 lk2=3.825626861e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.886133968e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.336345769e-8 nfactor=3.272300222e+00 lnfactor=-8.991423180e-7 eta0=1.556200358e-01 leta0=-1.494354750e-7 etab=-5.596804500e-02 letab=-2.772905143e-8 u0=3.355601231e-02 lu0=-8.171939531e-9 ua=-1.258399038e-10 lua=-1.322498677e-15 ub=8.990623895e-19 lub=1.318888206e-24 uc=5.360287210e-11 luc=2.076351371e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.430964044e+04 lvsat=-8.516435621e-3 a0=2.109817335e+00 la0=-1.135583262e-6 ags=1.494697789e-01 lags=9.971270444e-7 a1=0.0 a2=0.42385546 b0=4.164311393e-24 lb0=-4.064934266e-30 b1=0.0 keta=5.085943942e-02 lketa=-9.973614859e-08 wketa=-2.775557562e-23 pketa=3.122502257e-29 dwg=0.0 dwb=0.0 pclm=1.280914582e-01 lpclm=7.429649702e-7 pdiblc1=1.649323322e-01 lpdiblc1=4.447643207e-7 pdiblc2=6.380373791e-03 lpdiblc2=-3.026395354e-09 wpdiblc2=1.387778781e-23 pdiblcb=-4.921630060e-02 lpdiblcb=4.785470340e-8 drout=8.528408000e-01 ldrout=-5.786932471e-7 pscbe1=1.154740475e+09 lpscbe1=-7.174936905e+02 wpscbe1=-1.907348633e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.887283200e-09 lalpha0=5.555455173e-14 alpha1=6.342739440e-01 lalpha1=4.263040254e-7 beta0=1.320696502e+01 lbeta0=1.290485941e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.876870551e-01 lkt1=1.295694180e-7 kt2=-4.725934087e-02 lkt2=1.115524596e-8 at=1.633894479e+05 lat=-9.542651645e-2 ute=-1.987865646e+00 lute=7.949316238e-7 ua1=-5.141762198e-10 lua1=2.097147098e-15 pua1=1.654361225e-36 ub1=6.086990610e-19 lub1=-2.008681104e-24 uc1=1.034951732e-10 luc1=-1.158560798e-16 wuc1=1.033975766e-31 puc1=1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.41 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.728351421e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.687738636e-10 k1=4.392858589e-01 lk1=6.565994532e-8 k2=-6.791127560e-04 lk2=-1.917957525e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.934635650e-01 ldsub=6.494860950e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.283898860e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-5.255500608e-9 nfactor=1.921323762e+00 lnfactor=4.195944397e-7 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=-7.632783294e-23 peta0=2.879640970e-28 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.762200157e-02 lu0=-2.379538021e-9 ua=-1.371839134e-09 lua=-1.062339720e-16 ub=2.298097091e-18 lub=-4.675993133e-26 uc=7.398743477e-11 luc=8.654082393e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.721405808e+04 lvsat=4.721661776e-2 a0=4.193627844e-01 la0=5.145302813e-7 ags=1.158188796e+00 lags=1.248009777e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.631044528e-02 lketa=1.463759397e-8 dwg=0.0 dwb=0.0 pclm=1.355090508e+00 lpclm=-4.547529740e-7 pdiblc1=7.353854155e-01 lpdiblc1=-1.120754702e-7 pdiblc2=5.362028211e-03 lpdiblc2=-2.032351573e-9 pdiblcb=2.343260119e-02 lpdiblcb=-2.306050500e-08 wpdiblcb=1.387778781e-23 ppdiblcb=7.806255642e-30 drout=-4.446812800e-01 ldrout=6.878647659e-07 pdrout=4.440892099e-28 pscbe1=5.756251585e+07 lpscbe1=3.535012140e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.970567686e-06 lalpha0=2.957074856e-12 walpha0=-1.058791184e-27 palpha0=7.411538288e-34 alpha1=1.281452112e+00 lalpha1=-2.054298828e-7 beta0=1.120652299e+01 lbeta0=3.243189417e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.318729451e-01 lkt1=-2.252634408e-8 kt2=-3.479216166e-02 lkt2=-1.014416479e-9 at=8.375791069e+04 lat=-1.769530623e-2 ute=-1.097743715e+00 lute=-7.394843689e-8 ua1=2.198525948e-09 lua1=-5.508191447e-16 ub1=-2.277567454e-18 lub1=8.087075466e-25 uc1=-7.921055025e-11 luc1=6.248955431e-17 puc1=-2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.42 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.153678631e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.928258575e-8 k1=3.947279698e-01 lk1=8.687556041e-8 k2=4.280392337e-03 lk2=-2.154097416e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.095184973e-01 ldsub=1.049178783e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.343419918e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.421488753e-9 nfactor=2.600316138e+00 lnfactor=9.630172565e-8 eta0=0.49 etab=-0.000625 u0=2.811425844e-02 lu0=-2.613919240e-09 wu0=5.551115123e-23 ua=-1.145591476e-09 lua=-2.139586271e-16 ub=1.978807687e-18 lub=1.052652480e-25 uc=7.706502979e-11 luc=-5.999455450e-19 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.045937246e+05 lvsat=1.037337287e-2 a0=1.5 ags=2.238075265e+00 lags=-5.016927259e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.163195547e-02 lketa=-1.874083449e-9 dwg=0.0 dwb=0.0 pclm=4.711604765e-01 lpclm=-3.388206463e-8 pdiblc1=8.117032664e-01 lpdiblc1=-1.484131464e-7 pdiblc2=-2.522103509e-04 lpdiblc2=6.407895190e-10 pdiblcb=1.559088000e-01 lpdiblcb=-8.613719240e-08 wpdiblcb=5.551115123e-23 ppdiblcb=4.163336342e-29 drout=1.0 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.185727360e-06 lalpha0=2.584115772e-14 alpha1=0.85 beta0=1.701486070e+01 lbeta0=4.776307318e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.089088954e-01 lkt1=1.415324515e-8 kt2=-5.484301818e-02 lkt2=8.532518139e-9 at=6.821312074e+04 lat=-1.029387212e-2 ute=-2.132730218e+00 lute=4.188458967e-7 ua1=-1.764351194e-10 lua1=5.799853180e-16 ub1=2.034441167e-19 lub1=-3.725913786e-25 pub1=3.851859889e-46 uc1=5.317860243e-11 luc1=-5.456872969e-19 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.43 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.976466525e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.788878209e-08 wvth0=-3.386786373e-08 pvth0=7.658743231e-15 k1=4.930134021e-01 lk1=6.464968589e-8 k2=1.163993855e-02 lk2=-2.320523251e-08 wk2=-2.485145702e-08 pk2=5.619809086e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.296581543e-01 ldsub=-5.793162321e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=1.286776183e-02 lcdscd=-1.688729789e-9 cit=0.0 voff='-5.687790480e-03+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.151483523e-8 nfactor=9.471475546e-01 lnfactor=4.701426564e-07 wnfactor=5.926820371e-06 pnfactor=-1.340267451e-12 eta0=1.581403714e+00 leta0=-2.468056702e-7 etab=9.611909611e-02 letab=-2.187732292e-08 wetab=4.163336342e-23 petab=-1.301042607e-29 u0=-2.033475499e-02 lu0=8.342146862e-09 wu0=2.042023116e-08 pu0=-4.617749394e-15 ua=-4.068051533e-09 lua=4.469148005e-16 wua=-8.573060992e-17 pua=1.938677720e-23 ub=2.368417726e-18 lub=1.716039230e-26 wub=1.998290978e-24 pub=-4.518855286e-31 uc=-1.503555767e-10 luc=5.082804073e-17 wuc=4.046784666e-16 puc=-9.151236971e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.796808285e+05 lvsat=-6.606524461e-03 wvsat=-1.430761614e-01 pvsat=3.235467083e-8 a0=1.5 ags=-2.725047683e+00 lags=6.206480450e-07 wags=1.554312234e-21 pags=1.526556659e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.801076620e-01 lketa=7.692881892e-08 wketa=4.109482272e-07 pketa=-9.293018831e-14 dwg=0.0 dwb=0.0 pclm=5.565153056e-01 lpclm=-5.318386426e-08 wpclm=2.735489883e-07 ppclm=-6.185927401e-14 pdiblc1=-2.942002886e-01 lpdiblc1=1.016714599e-7 pdiblc2=-1.041058628e-02 lpdiblc2=2.937964019e-9 pdiblcb=-4.964630236e-01 lpdiblcb=6.138756232e-8 drout=2.107836980e+00 ldrout=-2.505218234e-7 pscbe1=8.191380802e+08 lpscbe1=-4.327808912e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.059378171e-05 lalpha0=-1.649386622e-12 alpha1=0.85 beta0=3.041889995e+01 lbeta0=-2.553505086e-06 wbeta0=8.924926207e-07 pbeta0=-2.018247113e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.016961167e-02 lkt1=-4.887974151e-08 wkt1=-4.462463104e-07 pkt1=1.009123556e-13 kt2=9.136848570e-03 lkt2=-5.935633008e-9 at=-6.212976870e+04 lat=1.918134752e-2 ute=2.035842074e+00 lute=-5.238183671e-07 wute=1.776356839e-21 pute=2.220446049e-28 ua1=7.768720193e-09 lua1=-1.216700324e-15 ub1=-6.244158411e-18 lub1=1.085443667e-24 uc1=-1.643023312e-10 luc1=4.863458112e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.44 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.68e-06 wmax=2.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.549813986e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=1.518388111e-8 k1=0.90707349 k2=-1.369819840e-01 wk2=1.114158165e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.958257461e+00 wnfactor=-2.657154186e-6 eta0=0.00069413878 etab=-0.043998 u0=3.309396652e-02 wu0=-9.154943007e-9 ua=-1.205708445e-09 wua=3.843535568e-17 ub=2.478324425e-18 wub=-8.958879980e-25 uc=1.751813957e-10 wuc=-1.814283231e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.373682007e+05 wvsat=6.414492044e-2 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.125962559e-01 wketa=-1.842392267e-7 dwg=0.0 dwb=0.0 pclm=2.158900541e-01 wpclm=-1.226394245e-7 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.406453525e+01 wbeta0=-4.001286279e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.432283650e-01 wkt1=2.000643140e-7 kt2=-0.028878939 at=60720.487 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.45 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.113909651e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.123654579e-07 wvth0=1.079181985e-08 pvth0=3.030207044e-13 k1=4.509691655e-01 lk1=6.516985304e-06 wk1=1.459086540e-07 pk1=-1.029337177e-11 k2=7.432822160e-03 lk2=-2.520072388e-06 wk2=-5.467183935e-08 pk2=3.996884008e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017280520e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.476438112e-07 wvoff=-3.167969614e-09 pvoff=-4.733385448e-13 nfactor=2.855212708e+00 lnfactor=-1.474726349e-05 wnfactor=-2.340901143e-07 pnfactor=2.419930727e-11 eta0=0.08 etab=-0.07 u0=3.177503734e-02 lu0=1.123728339e-07 wu0=-4.431371950e-10 pu0=-2.054048841e-13 ua=-7.599440421e-10 lua=-1.379098595e-15 wua=5.407358511e-17 pua=2.979659036e-21 ub=1.640904249e-18 lub=8.142629409e-24 wub=-6.681844800e-26 pub=-1.521124663e-29 uc=-7.946279064e-11 luc=5.618322440e-15 wuc=1.966905152e-16 puc=-8.205075772e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.070406966e+00 la0=1.040847049e-05 wa0=4.456853816e-07 pa0=-1.443371509e-11 ags=2.925775589e-01 lags=6.497800980e-06 wags=1.703035714e-07 pags=-1.002887809e-11 a1=0.0 a2=0.42385546 b0=-9.676380820e-24 lb0=3.572977822e-28 wb0=1.497228208e-29 pb0=-4.985599081e-34 b1=0.0 keta=-5.251190380e-03 lketa=-2.467254744e-07 wketa=-1.747328776e-09 pketa=4.253233787e-13 dwg=0.0 dwb=0.0 pclm=5.115884910e-02 lpclm=6.466704889e-07 wpclm=3.937366444e-08 ppclm=-7.865336756e-13 pdiblc1=0.39 pdiblc2=6.519696279e-03 lpdiblc2=-1.208370063e-07 wpdiblc2=-5.143550334e-09 ppdiblc2=1.678569801e-13 pdiblcb=9.806954753e+00 lpdiblcb=-2.630310212e-04 wpdiblcb=-1.507186282e-05 ppdiblcb=3.288183938e-10 drout=0.56 pscbe1=2.884416584e+08 lpscbe1=1.194071452e+04 wpscbe1=6.240318100e+02 ppscbe1=-1.549496892e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.383284327e-01 lkt1=-9.410351868e-07 wkt1=1.949766955e-08 pkt1=1.869037761e-12 kt2=-4.794737592e-02 lkt2=-1.044018015e-06 wkt2=2.171738047e-09 pkt2=1.889995471e-12 at=140000.0 ute=-1.881602031e+00 lute=-2.725108706e-05 wute=-4.159446421e-08 pute=4.840571214e-11 ua1=7.209456077e-10 lua1=-6.695541727e-14 wua1=-7.850376991e-16 pua1=1.124900486e-19 ub1=-1.152844987e-18 lub1=4.443852500e-23 wub1=1.042056652e-24 pub1=-6.974468188e-29 uc1=-4.396503424e-12 luc1=2.680225168e-15 wuc1=3.581457136e-17 puc1=-4.461565845e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.46 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.057659805e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.596095488e-8 k1=7.772076985e-01 wk1=-3.693747708e-7 k2=-1.187213244e-01 wk2=1.454111000e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.933106932e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' wvoff=-2.686316997e-8 nfactor=2.116968661e+00 wnfactor=9.773207044e-7 eta0=0.08 etab=-0.07 u0=3.740039121e-02 wu0=-1.072565049e-8 ua=-8.289813472e-10 wua=2.032345157e-16 ub=2.048522089e-18 wub=-8.282893664e-25 uc=2.017889209e-10 wuc=-2.140533730e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.591452202e+00 wa0=-2.768625169e-7 ags=6.178557299e-01 wags=-3.317393706e-7 a1=0.0 a2=0.42385546 b0=8.209850140e-24 wb0=-9.985492947e-30 b1=0.0 keta=-1.760220133e-02 wketa=1.954424527e-8 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=4.706282143e-04 wpdiblc2=3.259324983e-9 pdiblcb=-3.360307483e+00 wpdiblcb=1.388697615e-6 drout=0.56 pscbe1=8.861906187e+08 wpscbe1=-1.516421704e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.854364012e-01 wkt1=1.130611976e-7 kt2=-1.002106372e-01 wkt2=9.678440342e-8 at=140000.0 ute=-3.245784127e+00 wute=2.381582478e-6 ua1=-2.630824588e-09 wua1=4.846183907e-15 ub1=1.071735633e-18 wub1=-2.449343380e-24 uc1=1.297748482e-10 wuc1=-1.875302159e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.47 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.888921102e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.345882845e-07 wvth0=4.066118842e-08 pvth0=-1.172510620e-13 k1=8.131687922e-01 lk1=-2.868305740e-07 wk1=-4.333493544e-07 pk1=5.102699796e-13 k2=-1.282182141e-01 lk2=7.574848383e-08 wk2=1.673107877e-07 pk2=-1.746748870e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.167790395e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.104268781e-08 wvoff=-4.270898453e-08 pvoff=1.263883720e-13 nfactor=1.772105277e+00 lnfactor=2.750677251e-06 wnfactor=1.431954477e-06 pnfactor=-3.626220803e-12 eta0=0.08 etab=-0.07 u0=3.606554055e-02 lu0=1.064695042e-08 wu0=-8.298456304e-09 pu0=-1.935963096e-14 ua=-1.111259757e-09 lua=2.251490986e-15 wua=5.916963713e-16 pua=-3.098424591e-21 ub=2.340001023e-18 lub=-2.324875619e-24 wub=-1.191553621e-24 pub=2.897445097e-30 uc=2.405632926e-10 luc=-3.092696615e-16 wuc=-2.607037344e-16 puc=3.720896274e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.763232061e+00 la0=-1.370139517e-06 wa0=-3.293159120e-07 pa0=4.183754130e-13 ags=5.683301264e-01 lags=3.950229486e-07 wags=-2.609861654e-07 pags=-5.643371872e-13 a1=0.0 a2=0.42385546 b0=1.637072031e-23 lb0=-6.509221038e-29 wb0=-1.991141244e-29 pb0=7.917048383e-35 b1=0.0 keta=-4.345760672e-03 lketa=-1.057351736e-07 wketa=-1.023337145e-08 pketa=2.375103206e-13 dwg=0.0 dwb=0.0 pclm=-1.918176595e-01 lpclm=2.196218356e-06 wpclm=-2.087113809e-07 ppclm=1.664710358e-12 pdiblc1=0.39 pdiblc2=-2.953831242e-03 lpdiblc2=2.731395435e-08 wpdiblc2=7.189557173e-09 ppdiblc2=-3.134806646e-14 pdiblcb=-6.675716521e+00 lpdiblcb=2.644415339e-05 wpdiblcb=2.769110261e-06 ppdiblcb=-1.101035900e-11 drout=0.56 pscbe1=8.142000026e+08 lpscbe1=5.742069444e+02 wpscbe1=-4.439193428e+01 ppscbe1=-8.554424690e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.803797996e-01 lkt1=-4.033214272e-08 wkt1=1.083980456e-07 pkt1=3.719393489e-14 kt2=-9.612799359e-02 lkt2=-3.256372064e-08 wkt2=9.189338339e-08 pkt2=3.901144094e-14 at=140000.0 ute=-2.769448426e+00 lute=-3.799318332e-06 wute=1.557758950e-06 pute=6.570928497e-12 ua1=-2.166142124e-09 lua1=-3.706370531e-15 wua1=4.157799275e-15 pua1=5.490649443e-21 ub1=7.656477753e-19 lub1=2.441398380e-24 wub1=-2.069546179e-24 pub1=-3.029314127e-30 uc1=1.009927653e-10 luc1=2.295698080e-16 wuc1=-1.599265696e-16 puc1=-2.201704368e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.48 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.741301717e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.043298405e-07 wvth0=-7.876374788e-08 pvth0=3.575987265e-13 k1=8.258033443e-01 lk1=-3.370672714e-07 wk1=-4.672133721e-07 pk1=6.449179195e-13 k2=-1.551818002e-01 lk2=1.829593694e-07 wk2=2.090119177e-07 pk2=-3.404842514e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.644934323e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.682431159e-07 wvoff=9.497281463e-08 pvoff=-4.210531862e-13 nfactor=8.994323591e-01 lnfactor=6.220543455e-06 wnfactor=3.022266488e-06 pnfactor=-9.949517640e-12 eta0=0.08 etab=-0.07 u0=3.981504366e-02 lu0=-4.261583913e-09 wu0=-1.285915037e-08 pu0=-1.225691090e-15 ua=-1.332158241e-09 lua=3.129813399e-15 wua=1.319414700e-15 pua=-5.991931634e-21 ub=2.992797430e-18 lub=-4.920482916e-24 wub=-2.639789771e-24 pub=8.655828991e-30 uc=2.316169767e-10 luc=-2.736978929e-16 wuc=-2.853571810e-16 puc=4.701150836e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=-1.170902345e-01 la0=6.106277652e-06 wa0=1.878978242e-06 pa0=-8.362102472e-12 ags=2.335679244e-01 lags=1.726082991e-06 wags=-6.867175038e-08 pags=-1.329005456e-12 a1=0.0 a2=0.42385546 b0=-8.111890208e-24 lb0=3.225397868e-29 wb0=9.866346046e-30 pb0=-3.922993370e-35 b1=0.0 keta=-8.830851688e-02 lketa=2.281121641e-07 wketa=1.416357780e-07 pketa=-3.663420716e-13 dwg=0.0 dwb=0.0 pclm=3.704547550e-01 lpclm=-3.945323313e-08 wpclm=1.691371210e-07 ppclm=1.623333279e-13 pdiblc1=0.39 pdiblc2=4.275440790e-03 lpdiblc2=-1.430614430e-09 wpdiblc2=-3.478297903e-09 ppdiblc2=1.106877615e-14 pdiblcb=-0.025 drout=0.56 pscbe1=1.147432962e+09 lpscbe1=-7.507726199e+02 wpscbe1=-5.550167553e+02 ppscbe1=1.174871265e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.710108522e-01 lkt1=-7.758435171e-08 wkt1=9.158004335e-08 pkt1=1.040645990e-13 kt2=-9.784205172e-02 lkt2=-2.574839239e-08 wkt2=9.022363930e-08 pkt2=4.565057053e-14 at=1.534436066e+05 lat=-5.345360828e-02 wat=1.825973975e-02 pat=-7.260320858e-8 ute=-2.510701879e+00 lute=-4.828129792e-06 wute=9.366382773e-07 pute=9.040588764e-12 ua1=2.066007674e-09 lua1=-2.053397370e-14 wua1=-3.332602741e-15 pua1=3.527350655e-20 ub1=-3.516702540e-18 lub1=1.946860563e-23 wub1=5.272617693e-24 pub1=-3.222275622e-29 uc1=5.638247705e-11 luc1=4.069463810e-16 wuc1=-7.647380863e-17 puc1=-5.519899639e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.49 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='3.966554615e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.463843233e-07 wvth0=1.584915602e-07 pvth0=-1.112500289e-13 k1=7.232444938e-01 lk1=-1.343970348e-07 wk1=-1.521605605e-07 pk1=2.233071647e-14 k2=-8.586935061e-02 lk2=4.598854250e-08 wk2=4.311641718e-08 pk2=-1.265218058e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-07 wdsub=8.881784197e-22 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.410724960e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.044574812e-07 wvoff=-1.521228292e-07 pvoff=6.724141104e-14 nfactor=4.589353468e+00 lnfactor=-1.071242486e-06 wnfactor=-2.155070521e-06 pnfactor=2.816044065e-13 eta0=1.556201771e-01 leta0=-1.494357543e-07 weta0=-2.312722238e-13 peta0=4.570253672e-19 etab=-5.596804500e-02 letab=-2.772905143e-8 u0=4.791401884e-02 lu0=-2.026626032e-08 wu0=-2.349374764e-08 pu0=1.978971941e-14 ua=2.195974806e-09 lua=-3.842257326e-15 wua=-3.799143616e-15 pua=4.123035722e-21 ub=-1.652587243e-18 lub=4.259428972e-24 wub=4.175218364e-24 pub=-4.811553926e-30 uc=9.755077482e-11 luc=-8.764844988e-18 wuc=-7.191116217e-17 puc=4.831672182e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.250579846e+05 lvsat=-8.904070550e-02 wvsat=-6.667578212e-02 pvsat=1.317604134e-7 a0=4.119496706e+00 la0=-2.265794318e-06 wa0=-3.288402181e-06 pa0=1.849344008e-12 ags=-3.651560575e-01 lags=2.909243006e-06 wags=8.420729928e-07 pags=-3.128760930e-12 a1=0.0 a2=0.42385546 b0=1.622378042e-23 lb0=-1.583661612e-29 wb0=-1.973269209e-29 pb0=1.926179113e-35 b1=0.0 keta=2.757168205e-01 lketa=-4.912514101e-07 wketa=-3.679300853e-07 pketa=6.406293751e-13 dwg=0.0 dwb=0.0 pclm=-7.433166066e-01 lpclm=2.161510450e-06 wpclm=1.425869331e-06 ppclm=-2.321140435e-12 pdiblc1=-6.318451294e-01 lpdiblc1=2.019304947e-06 wpdiblc1=1.303752619e-06 ppdiblc1=-2.576392485e-12 pdiblc2=1.095896664e-02 lpdiblc2=-1.463817048e-08 wpdiblc2=-7.491869069e-09 ppdiblc2=1.900013862e-14 pdiblcb=-1.882408497e-01 lpdiblcb=3.225861198e-07 wpdiblcb=2.274833673e-07 ppdiblcb=-4.495380715e-13 drout=1.240960114e+00 ldrout=-1.345669796e-06 wdrout=-6.350726477e-07 pdrout=1.254989922e-12 pscbe1=2.182036796e+09 lpscbe1=-2.795290502e+03 wpscbe1=-1.680946478e+03 ppscbe1=3.399861523e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-8.291676297e-08 lalpha0=2.231388803e-13 walpha0=1.387633343e-13 palpha0=-2.742152203e-19 alpha1=-4.229498316e-01 lalpha1=2.515521988e-06 walpha1=1.729916234e-06 palpha1=-3.418549747e-12 beta0=1.131583479e+01 lbeta0=5.027616468e-06 wbeta0=3.094422354e-06 pbeta0=-6.114999413e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-5.666636745e-01 lkt1=3.090522339e-07 wkt1=2.928562207e-07 pkt1=-2.936845010e-13 kt2=-1.852391368e-01 lkt2=1.469601338e-07 wkt2=2.257738565e-07 pkt2=-2.222150934e-13 at=2.424843300e+05 lat=-2.294101872e-01 wat=-1.294215318e-01 pat=2.192350687e-7 ute=-8.285966809e+00 lute=6.584579146e-06 wute=1.030546957e-05 pute=-9.473496027e-12 ua1=-1.914313411e-08 lua1=2.137817490e-14 wua1=3.048222847e-14 pua1=-3.154919874e-20 ub1=1.585972640e-17 lub1=-1.882185315e-23 wub1=-2.495498152e-23 pub1=2.751109078e-29 uc1=6.271597049e-10 luc1=-7.209870469e-16 wuc1=-8.568628472e-16 puc1=9.901649091e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.50 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.317985559e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.446628380e-08 wvth0=6.714742742e-08 pvth0=-2.208573255e-14 k1=5.557583055e-01 lk1=2.909226309e-08 wk1=-1.905817679e-07 pk1=5.983504023e-14 k2=-2.167394797e-02 lk2=-1.667490105e-08 wk2=3.435347095e-08 pk2=-4.098353299e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.479196217e-01 ldsub=1.094056921e-07 wdsub=7.452273465e-08 pdsub=-7.274432412e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-4.565762667e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.635747399e-08 wvoff=-1.353733068e-07 pvoff=5.089159921e-14 nfactor=5.042173106e+00 lnfactor=-1.513256035e-06 wnfactor=-5.106589607e-06 pnfactor=3.162688441e-12 eta0=-4.616718742e-01 leta0=4.531252395e-07 weta0=4.625444475e-13 peta0=-2.202340631e-19 etab=-1.632660008e-01 letab=7.700834592e-08 wetab=-1.410113851e-09 petab=1.376462894e-15 u0=2.985084338e-02 lu0=-2.634144481e-09 wu0=-3.647013737e-09 pu0=4.166079678e-16 ua=-1.576921233e-09 lua=-1.593976788e-16 wua=3.355721464e-16 pua=8.699081638e-23 ub=2.541609194e-18 lub=1.653228380e-25 wub=-3.984544719e-25 pub=-3.470272179e-31 uc=1.055135756e-10 luc=-1.653762153e-17 wuc=-5.158565684e-17 puc=2.847626436e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-5.918801558e+04 lvsat=9.080844816e-02 wvsat=1.413781579e-01 pvsat=-7.132852742e-8 a0=2.082381437e+00 la0=-2.772927679e-07 wa0=-2.721167487e-06 pa0=1.295645803e-12 ags=3.731744844e+00 lags=-1.089889452e-06 wags=-4.211063437e-06 pags=1.803787452e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-3.995377377e-01 lketa=1.678888733e-07 wketa=5.452538204e-07 pketa=-2.507623099e-13 dwg=0.0 dwb=0.0 pclm=2.766725258e+00 lpclm=-1.264767775e-06 wpclm=-2.309832532e-06 ppclm=1.325412638e-12 pdiblc1=1.342014350e+00 lpdiblc1=9.254964994e-08 wpdiblc1=-9.926160061e-07 ppdiblc1=-3.348244008e-13 pdiblc2=-7.510332783e-03 lpdiblc2=3.390377589e-09 wpdiblc2=2.106281259e-08 ppdiblc2=-8.873114118e-15 pdiblcb=3.014816994e-01 lpdiblcb=-1.554496904e-07 wpdiblcb=-4.549667345e-07 ppdiblcb=2.166260411e-13 drout=-1.220919908e+00 ldrout=1.057459922e-06 wdrout=1.270145295e-06 pdrout=-6.047619004e-13 pscbe1=-2.092469265e+09 lpscbe1=1.377208746e+03 wpscbe1=3.518058303e+03 ppscbe1=-1.675074208e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.165315590e-05 lalpha0=1.151726583e-11 walpha0=1.420716281e-11 palpha0=-1.400688641e-17 alpha1=3.395899663e+00 lalpha1=-1.212194482e-06 walpha1=-3.459832468e-06 palpha1=1.647350792e-12 beta0=3.522293653e+00 lbeta0=1.263517254e-05 wbeta0=1.257356615e-05 pbeta0=-1.536793292e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.990952945e-01 lkt1=-4.974449421e-08 wkt1=-5.363347965e-08 pkt1=4.453656913e-14 kt2=-3.097782830e-02 lkt2=-3.619882884e-09 wkt2=-6.241325025e-09 pkt2=4.263277779e-15 at=-2.004109801e+04 lat=2.685033402e-02 wat=1.698444496e-01 pat=-7.288922932e-8 ute=-1.739299944e+00 lute=1.941419392e-07 wute=1.049766909e-06 pute=-4.386714567e-13 ua1=4.535025217e-09 lua1=-1.734928828e-15 wua1=-3.823171697e-15 pua1=1.937537360e-21 ub1=-6.407326370e-18 lub1=2.913818675e-24 wub1=6.757450178e-24 pub1=-3.444555447e-30 uc1=-3.025200316e-10 luc1=1.865068124e-16 wuc1=3.653972848e-16 puc1=-2.029272071e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.51 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.989188996e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.749212820e-08 wvth0=2.691514276e-08 pvth0=-2.929693463e-15 k1=8.060266948e-01 lk1=-9.006952671e-08 wk1=-6.730007004e-07 pk1=2.895320610e-13 k2=-1.533906408e-01 lk2=4.604015822e-08 wk2=2.579942735e-07 pk2=-1.105817905e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.002345918e-01 ldsub=2.275608468e-07 wdsub=3.432152042e-07 pdsub=-2.006784818e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=-3.370010952e-03 lcdscd=4.175717935e-09 wcdscd=1.435021106e-08 pcdscd=-6.832652094e-15 cit=0.0 voff='-1.887515309e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.177468520e-08 wvoff=8.902934945e-08 pvoff=-5.595458391e-14 nfactor=-1.052028069e+00 lnfactor=1.388412535e-06 wnfactor=5.976265084e-06 pnfactor=-2.114257660e-12 eta0=-7.917257321e-01 leta0=6.102757632e-07 weta0=2.097264744e-06 peta0=-9.985832464e-13 etab=-1.159631597e-01 letab=5.448576041e-08 wetab=1.887257547e-07 petab=-8.915406901e-14 u0=5.344024449e-02 lu0=-1.386590757e-08 wu0=-4.144045510e-08 pu0=1.841142596e-14 ua=6.572337766e-10 lua=-1.223159308e-15 wua=-2.949930510e-15 pua=1.651336909e-21 ub=1.575914872e-18 lub=6.251246697e-25 wub=6.592462614e-25 pub=-8.506366142e-31 uc=1.150341124e-10 luc=-2.107069180e-17 wuc=-6.212812636e-17 puc=3.349591362e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.440334061e+05 lvsat=-5.952586690e-03 wvsat=-6.453444100e-02 pvsat=2.671387377e-8 a0=1.5 ags=5.953233758e+00 lags=-2.147620298e-06 wags=-6.079046970e-06 pags=2.693201659e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.665092979e-01 lketa=5.693564410e-08 wketa=2.206973675e-07 pketa=-9.622929862e-14 dwg=0.0 dwb=0.0 pclm=-2.971661992e-01 lpclm=1.940612477e-07 wpclm=1.257199110e-06 ppclm=-3.729795390e-13 pdiblc1=3.313561455e+00 lpdiblc1=-8.461749024e-07 wpdiblc1=-4.093745520e-06 ppdiblc1=1.141735002e-12 pdiblc2=1.218033609e-02 lpdiblc2=-5.985058727e-09 wpdiblc2=-2.034315196e-08 ppdiblc2=1.084175622e-14 pdiblcb=4.747103024e-01 lpdiblcb=-2.379300645e-07 wpdiblcb=-5.216491600e-07 ppdiblcb=2.483759444e-13 drout=-3.010246809e-01 ldrout=6.194646874e-07 wdrout=2.128843267e-06 pdrout=-1.013618918e-12 pscbe1=7.775245680e+08 lpscbe1=1.070136230e+01 wpscbe1=3.677614484e+01 ppscbe1=-1.751044650e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.230242466e-05 lalpha0=1.111515241e-13 walpha0=-1.491748770e-11 palpha0=-1.395918170e-19 alpha1=0.85 beta0=2.735601155e+01 lbeta0=1.287081431e-06 wbeta0=-1.692103899e-05 pbeta0=-1.324489608e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.413124179e-01 lkt1=1.797019807e-08 wkt1=5.302130068e-08 pkt1=-6.245611361e-15 kt2=-8.882559683e-02 lkt2=2.392352224e-08 wkt2=5.560508177e-08 pkt2=-2.518402296e-14 at=6.449632294e+04 lat=-1.340097544e-02 wat=6.081729330e-03 pat=5.084097239e-9 ute=-5.002565161e+00 lute=1.747899986e-06 wute=4.695859259e-06 pute=-2.174707284e-12 ua1=-6.781547933e-09 lua1=3.653299046e-15 wua1=1.080782720e-14 pua1=-5.028807933e-21 ub1=6.395571014e-18 lub1=-3.182101674e-24 wub1=-1.013206578e-23 pub1=4.597151125e-30 uc1=3.765168716e-10 luc1=-1.368071026e-16 wuc1=-5.290725897e-16 puc1=2.229621011e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.52 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.861294744e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.721357874e-08 wvth0=-1.502251251e-08 pvth0=6.553920151e-15 k1=-7.060671499e-01 lk1=2.518693270e-07 wk1=1.962033924e-06 pk1=-3.063441287e-13 k2=4.775180688e-01 lk2=-9.663101375e-08 wk2=-7.871594558e-07 pk2=1.257650933e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.904090211e+00 ldsub=-2.256891467e-07 wdsub=-1.758073834e-06 pdsub=2.744986161e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=4.418922952e-02 lcdscd=-6.579138468e-09 wcdscd=-5.125075379e-08 pcdscd=8.002087694e-15 cit=0.0 voff='3.070581870e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.034574117e-08 wvoff=-5.117406135e-07 pvoff=7.990113243e-14 nfactor=1.159930070e+01 lnfactor=-1.472508348e-06 wnfactor=-1.150310609e-05 pnfactor=1.838457420e-12 eta0=6.158995614e+00 leta0=-9.615325591e-07 weta0=-7.490231230e-06 peta0=1.169494743e-12 etab=5.018855292e-01 letab=-8.523207072e-08 wetab=-6.639483107e-07 petab=1.036662334e-13 u0=-9.189377640e-02 lu0=1.899934658e-08 wu0=1.375109698e-07 pu0=-2.205593346e-14 ua=-1.269058834e-08 lua=1.795263794e-15 wua=1.402317116e-14 pua=-2.186892410e-21 ub=1.059986038e-17 lub=-1.415514271e-24 wub=-1.147067046e-23 pub=1.892374234e-30 uc=3.517486663e-11 luc=-3.011641408e-18 wuc=1.010983416e-16 puc=-3.415466940e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.135073598e+04 lvsat=2.918536167e-02 wvsat=1.695053490e-01 pvsat=-2.621094819e-8 a0=1.5 ags=-1.423642612e+01 lags=2.417988629e-06 wags=1.883586134e-05 pags=-2.940956046e-12 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.754556789e-01 lketa=-4.300854788e-08 wketa=-6.617382673e-07 pketa=1.033211661e-13 dwg=0.0 dwb=0.0 pclm=1.497935204e+00 lpclm=-2.118758031e-07 wpclm=-1.266879446e-06 ppclm=1.978054891e-13 pdiblc1=-2.179936755e+00 lpdiblc1=3.961028088e-07 wpdiblc1=3.085596637e-06 ppdiblc1=-4.817727165e-13 pdiblc2=-6.490204233e-02 lpdiblc2=1.144604200e-08 wpdiblc2=8.916338869e-08 ppdiblc2=-1.392161486e-14 pdiblcb=-1.635039818e+00 lpdiblcb=2.391603887e-07 wpdiblcb=1.863032714e-06 ppdiblcb=-2.908864758e-13 drout=6.754353698e+00 ldrout=-9.760103575e-07 wdrout=-7.603011667e-06 pdrout=1.187103830e-12 pscbe1=8.994074803e+08 lpscbe1=-1.686075196e+01 wpscbe1=-1.313433744e+02 ppscbe1=2.050742911e-5 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=4.126412212e-05 lalpha0=-6.438130891e-12 walpha0=-5.018532593e-11 palpha0=7.835736050e-18 alpha1=0.85 beta0=7.612893730e+01 lbeta0=-9.742232906e-06 wbeta0=-7.390201872e-05 pbeta0=1.156096122e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.530414395e-01 lkt1=2.062255210e-08 wkt1=8.206304986e-08 pkt1=-1.281299635e-14 kt2=1.192271299e-01 lkt2=-2.312468917e-08 wkt2=-1.801387456e-07 pkt2=2.812614319e-14 at=-2.477114787e+05 lat=5.720044798e-02 wat=3.036640115e-01 pat=-6.220996973e-8 ute=1.175128629e+01 lute=-2.040748965e-06 wute=-1.589720649e-05 pute=2.482126233e-12 ua1=3.033529071e-08 lua1=-4.740154379e-15 wua1=-3.692527315e-14 pua1=5.765364448e-21 ub1=-2.637626537e-17 lub1=4.228790318e-24 wub1=3.294180424e-23 pub1=-5.143401546e-30 uc1=-1.066345080e-09 luc1=1.894759278e-16 wuc1=1.475996313e-15 puc1=-2.304561604e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.53 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.26e-06 wmax=1.68e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.477886770e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' wvth0=2.695320193e-8 k1=0.90707349 k2=-1.413719613e-01 wk2=1.832482244e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.168366466e+00 wnfactor=2.716122316e-7 eta0=0.00069413878 etab=-0.043998 u0=2.979082280e-02 wu0=-3.750068390e-9 ua=-1.192511062e-09 wua=1.684071653e-17 ub=1.533954559e-18 wub=6.493674149e-25 uc=1.588628867e-11 wuc=7.922339325e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.755719575e+05 wvsat=1.632800816e-3 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=0.0 dwg=0.0 dwb=0.0 pclm=0.14094 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=1.373312271e+01 wbeta0=1.421557388e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=1.186386775e+05 wat=-9.477049255e-2 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.54 nmos lmin=2.0e-05 lmax=0.0001 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.707480052e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.869322339e-06 wvth0=-1.830312796e-07 pvth0=3.656257733e-12 k1=4.949059275e-01 lk1=-4.272885007e-07 wk1=9.246916123e-08 pk1=-1.847176541e-12 k2=-7.087086284e-03 lk2=1.582016719e-07 wk2=-3.701153607e-08 pk2=7.393474782e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.270573901e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.737860854e-07 wvoff=-1.414164645e-08 pvoff=2.824954527e-13 nfactor=-2.378170621e-01 lnfactor=6.309097116e-05 wnfactor=3.527906321e-06 pnfactor=-7.047393646e-11 eta0=0.08 etab=-0.07 u0=6.121108038e-02 lu0=-6.518029472e-07 wu0=-3.624566649e-08 pu0=7.240483633e-13 ua=8.888569869e-10 lua=-3.097786180e-14 wua=-1.951333428e-15 pua=3.898010194e-20 ub=1.336014698e-18 lub=6.293741821e-25 wub=3.040132251e-25 pub=-6.073009531e-30 uc=1.853722886e-10 luc=-3.187657714e-15 wuc=-1.254236246e-16 puc=2.505479383e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.711015575e+00 la0=-6.935586063e-06 wa0=-3.334753380e-07 pa0=6.661548704e-12 ags=7.554309923e-01 lags=-8.196687873e-06 wags=-3.926567282e-07 pags=7.843764204e-12 a1=0.0 a2=0.42385546 b0=-1.072251100e-07 lb0=2.141943380e-12 wb0=1.304159712e-13 pb0=-2.605207178e-18 b1=-1.797840772e-08 lb1=3.591391176e-13 wb1=2.186681370e-14 pb1=-4.368144443e-19 keta=-1.179579840e-02 lketa=2.050039111e-07 wketa=6.212760153e-09 pketa=-1.241069417e-13 dwg=0.0 dwb=0.0 pclm=3.899094693e-01 lpclm=-6.120257970e-06 wpclm=-3.726426174e-07 ppclm=7.443959605e-12 pdiblc1=0.39 pdiblc2=9.195559666e-03 lpdiblc2=-1.207594770e-07 wpdiblc2=-8.398154805e-09 ppdiblc2=1.677626825e-13 pdiblcb=-1.401431107e+01 lpdiblcb=2.356337033e-04 wpdiblcb=1.390151402e-05 ppdiblcb=-2.776985346e-10 drout=0.56 pscbe1=3.414639747e+09 lpscbe1=-5.299920474e+04 wpscbe1=-3.178306654e+03 ppscbe1=6.349028596e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.600064000e-01 lkt1=3.346530151e-06 wkt1=1.674923910e-07 pkt1=-3.345850783e-12 kt2=-9.922157029e-02 lkt2=1.569822975e-06 wkt2=6.453561772e-08 pkt2=-1.289172276e-12 at=-2.087443630e+04 lat=3.213649618e+00 wat=1.956686811e-01 pat=-3.908704185e-6 ute=-5.017918848e+00 lute=7.451535901e-05 wute=3.773051226e-06 pute=-7.537098442e-11 ua1=-3.556212340e-09 lua1=9.807907904e-14 wua1=4.417192524e-15 pua1=-8.823843859e-20 ub1=3.672190917e-19 lub1=-2.615433720e-23 wub1=-8.067699250e-25 pub1=1.611614574e-29 uc1=-6.067838646e-11 luc1=7.245357204e-16 wuc1=1.042692126e-16 puc1=-2.082895972e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.55 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.5271105+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.47351598 k2=0.0008324469 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.11141737+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=2.9205 eta0=0.08 etab=-0.07 u0=0.028582 ua=-6.6188645e-10 ub=1.367521e-18 uc=2.5799e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.363822 ags=0.345107 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.0015333577 dwg=0.0 dwb=0.0 pclm=0.083531 pdiblc1=0.39 pdiblc2=0.0031503727 pdiblcb=-2.2185512 drout=0.56 pscbe1=761513800.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.29248 kt2=-0.020636654 at=140000.0 ute=-1.2877 ua1=1.3536e-9 ub1=-9.4206e-19 uc1=-2.4408323e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.56 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.223228346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.818707001e-8 k1=4.568785944e-01 lk1=1.327020504e-7 k2=9.340993149e-03 lk2=-6.786532205e-08 wk2=-1.734723476e-24 pk2=6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.167922808e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.287101972e-08 wvoff=-1.110223025e-22 nfactor=2.949426389e+00 lnfactor=-2.307208158e-7 eta0=0.08 etab=-0.07 u0=2.924273440e-02 lu0=-5.270107433e-9 ua=-6.247801648e-10 lua=-2.959647776e-16 ub=1.360332146e-18 lub=5.733927629e-26 uc=2.621848235e-11 luc=-3.345848257e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.492475844e+00 la0=-1.026160561e-6 ags=3.537531077e-01 lags=-6.896253114e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.275941100e-02 lketa=8.954052784e-08 wketa=-1.734723476e-24 pketa=1.387778781e-29 dwg=0.0 dwb=0.0 pclm=-3.634155134e-01 lpclm=3.564906175e-06 wpclm=1.110223025e-22 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=2.957262709e-03 lpdiblc2=1.540271552e-9 pdiblcb=-4.399015674e+00 lpdiblcb=1.739168118e-5 drout=0.56 pscbe1=7.777019419e+08 lpscbe1=-1.291188214e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912573382e-01 lkt1=-9.752116958e-9 kt2=-2.057529825e-02 lkt2=-4.893818432e-10 at=140000.0 ute=-1.488693675e+00 lute=1.603152885e-6 ua1=1.252307935e-09 lua1=8.079192830e-16 ub1=-9.358870489e-19 lub1=-4.923629781e-26 uc1=-3.049530213e-11 luc1=4.855057335e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.57 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.093723706e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.967987643e-8 k1=4.416709045e-01 lk1=1.931698936e-7 k2=1.666314832e-02 lk2=-9.697920683e-08 pk2=-2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.640889714e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.793744597e-8 nfactor=3.384272625e+00 lnfactor=-1.959728587e-6 eta0=0.08 etab=-0.07 u0=2.924253632e-02 lu0=-5.269319858e-09 wu0=-2.775557562e-23 ua=-2.473648295e-10 lua=-1.796619479e-15 ub=8.224210119e-19 lub=2.196147102e-24 uc=-2.997348756e-12 luc=1.128202696e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.427763872e+00 la0=-7.688569563e-7 ags=1.771075391e-01 lags=6.334042736e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.814126858e-02 lketa=-7.308613666e-08 wketa=1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.095155328e-01 lpclm=9.401361739e-8 pdiblc1=0.39 pdiblc2=1.415661641e-03 lpdiblc2=7.669887058e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.911105335e+08 lpscbe1=2.151803947e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.957157780e-01 lkt1=7.975246273e-9 kt2=-2.366218282e-02 lkt2=1.178449104e-8 at=1.684563584e+05 lat=-1.131463511e-1 ute=-1.740618726e+00 lute=2.604841151e-6 ua1=-6.739841536e-10 lua1=8.467118605e-15 ub1=8.183264192e-19 lub1=-7.024227620e-24 pub1=3.081487911e-45 uc1=-6.492586981e-12 luc1=-4.688748644e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.58 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.269636961e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.491702467e-8 k1=5.981414663e-01 lk1=-1.160372166e-7 k2=-5.041999168e-02 lk2=3.558620112e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.009647561e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.917308910e-8 nfactor=2.817502433e+00 lnfactor=-8.397136079e-7 eta0=1.556199869e-01 leta0=-1.494353785e-7 etab=-5.596804500e-02 letab=-2.772905143e-8 u0=2.859798223e-02 lu0=-3.995593312e-9 ua=-9.275965507e-10 lua=-4.523890865e-16 ub=1.780184404e-18 lub=3.034763837e-25 uc=3.842701720e-11 luc=3.096008872e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.023864000e+04 lvsat=1.928977490e-2 a0=1.415845595e+00 la0=-7.453048199e-7 ags=3.271776224e-01 lags=3.368453795e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.678710971e-02 lketa=3.545980911e-08 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=4.290014341e-01 lpclm=2.531204263e-7 pdiblc1=4.400712671e-01 lpdiblc1=-9.894763339e-8 pdiblc2=4.799318577e-03 lpdiblc2=9.833207738e-10 pdiblcb=-1.209086295e-03 lpdiblcb=-4.701408105e-8 drout=7.188175127e-01 ldrout=-3.138450042e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.117136320e-08 lalpha0=-2.314772989e-15 alpha1=9.993488080e-01 lalpha1=-2.951335560e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.258838054e-01 lkt1=6.759137127e-8 kt2=3.871048534e-04 lkt2=-3.574017210e-8 at=1.360768260e+05 lat=-4.915999135e-02 wat=-1.164153218e-16 ute=1.869609889e-01 lute=-1.204318517e-6 ua1=5.918675958e-09 lua1=-4.560874379e-15 ub1=-4.657704193e-18 lub1=3.797153610e-24 uc1=-7.733386419e-11 luc1=9.310451173e-17 wuc1=-5.169878828e-32 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.59 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.870056768e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.692114131e-9 k1=3.990662161e-01 lk1=7.828730192e-8 k2=6.570711535e-03 lk2=-2.004447595e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.091905561e-01 ldsub=4.959692731e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.569585476e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.484466620e-9 nfactor=8.436487450e-01 lnfactor=1.087036036e-6 eta0=-4.616714939e-01 leta0=4.531250584e-07 weta0=4.510281038e-23 peta0=8.153200337e-29 etab=-1.644253650e-01 letab=7.814004309e-8 u0=2.685234983e-02 lu0=-2.291618679e-9 ua=-1.301021280e-09 lua=-8.787576494e-17 ub=2.214008792e-18 lub=-1.199952198e-25 uc=6.310099629e-11 luc=6.874929471e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.704996039e+04 lvsat=3.216371986e-2 a0=-1.549019290e-01 la0=7.879583848e-7 ags=2.695021758e-01 lags=3.931444592e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.875782245e-02 lketa=-3.828231879e-08 wketa=-1.387778781e-23 pketa=6.938893904e-30 dwg=0.0 dwb=0.0 pclm=8.676323403e-01 lpclm=-1.750429920e-7 pdiblc1=5.259075539e-01 lpdiblc1=-1.827355231e-07 wpdiblc1=-4.440892099e-22 pdiblc2=9.807043116e-03 lpdiblc2=-3.904899426e-9 pdiblcb=-7.258182741e-02 lpdiblcb=2.265542098e-8 drout=-1.766347053e-01 ldrout=5.602381421e-07 pdrout=2.220446049e-28 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.765727360e-08 lalpha0=1.115456377e-15 alpha1=5.513023840e-01 lalpha1=1.422206881e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.431915482e-01 lkt1=-1.312751794e-8 kt2=-3.610930687e-02 lkt2=-1.147107452e-10 at=1.196012296e+05 lat=-3.307756865e-2 ute=-8.762049469e-01 lute=-1.665239728e-7 ua1=1.391698507e-09 lua1=-1.419287174e-16 ub1=-8.515011762e-19 lub1=8.178182225e-26 wub1=7.703719778e-40 uc1=-2.098513587e-12 luc1=1.966457754e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.60 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.210479312e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.990085699e-8 k1=2.527004922e-01 lk1=1.479772922e-7 k2=5.872651086e-02 lk2=-4.487772962e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.819493130e-01 ldsub=6.256746383e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413312e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.155535806e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.422992879e-8 nfactor=3.861524120e+00 lnfactor=-3.498830736e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.920295691e-02 letab=-1.881473159e-08 wetab=-9.540979118e-24 petab=-3.144186300e-30 u0=1.936882429e-02 lu0=1.271557234e-9 ua=-1.768133457e-09 lua=1.345331586e-16 wua=-1.654361225e-30 ub=2.117932481e-18 lub=-7.424982916e-26 uc=6.395374912e-11 luc=6.468903149e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.097462453e+04 lvsat=1.601096598e-2 a0=1.5 ags=9.551765888e-01 lags=6.667018692e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.494316756e-02 lketa=-2.218194427e-8 dwg=0.0 dwb=0.0 pclm=7.364749379e-01 lpclm=-1.125942310e-7 pdiblc1=-5.222503249e-02 lpdiblc1=9.253421406e-8 pdiblc2=-4.545350845e-03 lpdiblc2=2.928792025e-09 wpdiblc2=1.734723476e-24 ppdiblc2=-8.673617380e-31 pdiblcb=4.582196898e-02 lpdiblcb=-3.372088902e-8 drout=1.449262890e+00 ldrout=-2.139102352e-7 pscbe1=8.077610961e+08 lpscbe1=-3.695337236e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.759816960e-08 lalpha0=-3.617762081e-15 alpha1=0.85 beta0=1.344390976e+01 lbeta0=1.981155425e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.977194842e-01 lkt1=1.283519537e-8 kt2=-4.310833573e-02 lkt2=3.217778860e-9 at=6.949658549e+04 lat=-9.220943808e-3 ute=-1.141734153e+00 lute=-4.009595862e-8 ua1=2.104407137e-09 lua1=-4.812749535e-16 ub1=-1.934788051e-18 lub1=5.975737015e-25 wub1=-7.703719778e-40 pub1=1.925929944e-46 uc1=-5.847484063e-11 luc1=4.650737639e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.61 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='8.823857636e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-7.899874906e-08 wvth0=-2.537255045e-07 pvth0=5.737647068e-14 k1=0.90707349 k2=-2.164108118e-01 lk2=1.734072397e-08 wk2=5.685375095e-08 pk2=-1.285667983e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586410187e-01 ldsub=-2.491733918e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.136835600e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280776e-8 nfactor=-7.036451375e+00 lnfactor=2.114541513e-06 wnfactor=1.116322372e-05 pnfactor=-2.524406760e-12 eta0=6.941427212e-04 leta0=-6.153674857e-16 etab=-0.043998 u0=1.748935937e-02 lu0=1.696571914e-09 wu0=4.470230690e-09 pu0=-1.010880087e-15 ua=-1.154436704e-09 lua=-4.245770439e-18 wua=-8.042423965e-18 pua=1.818681586e-24 ub=6.649713698e-20 lub=3.896535538e-25 wub=1.340869643e-24 pub=-3.032188976e-31 uc=3.575855327e-10 luc=-5.993181387e-17 wuc=-2.910439482e-16 puc=6.581551426e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.385382466e+05 lvsat=5.255118741e-03 wvsat=-1.280192249e-02 pvsat=2.894975543e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.885609012e-01 lketa=1.142920518e-07 wketa=3.891495467e-07 pketa=-8.800072189e-14 dwg=0.0 dwb=0.0 pclm=3.637956964e-01 lpclm=-2.831803807e-08 wpclm=1.125540227e-07 ppclm=-2.545251649e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-6.604864909e-08 lalpha0=1.982051491e-14 walpha0=8.381682544e-14 palpha0=-1.895400164e-20 alpha1=0.85 beta0=1.725522692e+01 lbeta0=-6.637604737e-07 wbeta0=-2.294984506e-06 pbeta0=5.189786163e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.496479997e-01 lkt1=4.719170217e-08 wkt1=1.995638701e-07 pkt1=-4.512857533e-14 kt2=-0.028878939 at=1.660312896e+05 lat=-3.105091565e-02 wat=-1.995638701e-01 pat=4.512857533e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.62 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=1.0e-06 wmax=1.26e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='3.188143043e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.379559551e-08 wvth0=5.328136997e-07 pvth0=-6.543061450e-14 k1=0.90707349 k2=-5.039519017e-02 lk2=-8.580291123e-09 wk2=-9.232858671e-08 pk2=1.043605365e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45862506 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.118353774e+01 lnfactor=-3.852974707e-06 wnfactor=-3.501901831e-05 pnfactor=4.686303782e-12 eta0=0.00069413878 etab=-0.043998 u0=2.879608017e-02 lu0=-6.881424387e-11 wu0=-2.540180833e-09 pu0=8.369752616e-17 ua=-1.178876828e-09 lua=-4.297872073e-19 wua=2.576422700e-19 pua=5.227424441e-25 ub=1.121291289e-18 lub=2.249622141e-25 wub=1.151282322e-24 pub=-2.736174917e-31 uc=-4.773210041e-10 luc=7.042715317e-17 wuc=6.791025457e-16 puc=-8.565927871e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.151987049e+05 lvsat=-6.714338574e-03 wvsat=-4.656449874e-02 pvsat=8.166529149e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=7.465502318e-01 lketa=-9.416686003e-08 wketa=-9.080156090e-07 pketa=1.145334569e-13 dwg=0.0 dwb=0.0 pclm=1.824279268e-01 wpclm=-5.046101855e-8 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.907954345e-07 lalpha0=-2.028209293e-14 walpha0=-1.955725927e-13 palpha0=2.466874455e-20 alpha1=0.85 beta0=9.447267864e+00 lbeta0=5.553430207e-07 wbeta0=5.354963848e-06 pbeta0=-6.754537199e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=1.618855327e-01 lkt1=-4.829069745e-08 wkt1=-4.656490302e-07 pkt1=5.873510608e-14 kt2=-0.028878939 at=-3.421257857e+05 lat=4.829069745e-02 wat=4.656490302e-01 pat=-5.873510608e-8 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.63 nmos lmin=2.0e-05 lmax=0.0001 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.318551619e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.702352679e-06 wvth0=4.541764642e-08 pvth0=-4.540680796e-12 k1=7.090279257e-01 lk1=-1.409865527e-05 wk1=-1.122918515e-07 pk1=1.122650541e-11 k2=-9.215278855e-02 lk2=5.566455559e-06 wk2=4.433526382e-08 pk2=-4.432468365e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.035923811e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.684340787e-07 wvoff=-3.730946603e-09 pvoff=3.730056250e-13 nfactor=3.979274815e+00 lnfactor=-6.338235233e-05 wnfactor=-5.048227337e-07 pnfactor=5.047022628e-11 eta0=0.08 etab=-0.07 u0=1.806428851e-02 lu0=6.296308583e-07 wu0=5.014833931e-09 pu0=-5.013637191e-13 ua=-1.638741430e-09 lua=5.847831441e-14 wua=4.657634413e-16 pua=-4.656522915e-20 ub=1.938728517e-18 lub=-3.419468956e-23 wub=-2.723511518e-25 pub=2.722861579e-29 uc=8.247136757e-11 luc=-3.392626948e-15 wuc=-2.702132608e-17 puc=2.701487771e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.360776278e+00 la0=1.823287066e-07 wa0=1.452197224e-09 pa0=-1.451850671e-13 ags=3.445412234e-01 lags=3.386957151e-08 wags=2.697616774e-10 pags=-2.696973014e-14 a1=0.0 a2=0.42385546 b0=5.814288815e-08 lb0=-3.480657992e-12 wb0=-2.772246877e-14 pb0=2.771585308e-18 b1=9.748803700e-09 lb1=-5.836010662e-13 wb1=-4.648219493e-15 pb1=4.647110242e-19 keta=-9.043586181e-03 lketa=4.495913021e-07 wketa=3.580869151e-09 pketa=-3.580014612e-13 dwg=0.0 dwb=0.0 pclm=-8.260293143e-02 lpclm=9.945419202e-06 wpclm=7.921248620e-08 ppclm=-7.919358293e-12 pdiblc1=0.39 pdiblc2=-2.308113044e-03 lpdiblc2=3.267660523e-07 wpdiblc2=2.602600341e-09 ppdiblc2=-2.601979257e-13 pdiblcb=3.248672826e+00 lpdiblcb=-3.272891596e-04 wpdiblcb=-2.606766745e-06 ppdiblcb=2.606144666e-10 drout=0.56 pscbe1=-5.756973567e+08 lpscbe1=8.005062783e+04 wpscbe1=6.375808926e+02 ppscbe1=-6.374287403e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.772763127e-01 lkt1=-9.101514812e-07 wkt1=-7.249102343e-09 pkt1=7.247372418e-13 kt2=-4.277241768e-02 lkt2=1.325132363e-06 wkt2=1.055430917e-08 pkt2=-1.055179049e-12 at=2.272342715e+05 lat=-5.222180630e+00 wat=-4.159321017e-02 pat=4.158328436e-6 ute=-8.582581435e-01 lute=-2.570804922e-05 wute=-2.047574318e-07 pute=2.047085685e-11 ua1=7.738659558e-10 lua1=3.470512042e-14 wua1=2.764165910e-16 pua1=-2.763506269e-20 ub1=-1.341379391e-20 lub1=-5.559235088e-23 wub1=-4.427775479e-25 pub1=4.426718835e-29 uc1=1.207163183e-10 luc1=-8.687721902e-15 wuc1=-6.919527847e-17 puc1=6.917876571e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.64 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='8.437370908e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.525456749e-06 wvth0=-3.027843095e-07 pvth0=2.415048831e-12 k1=-3.093204041e-01 lk1=6.244009465e-06 wk1=7.486123430e-07 pk1=-5.971033859e-12 k2=3.099132677e-01 lk2=-2.465270662e-06 wk2=-2.955684255e-07 pk2=2.357493959e-12 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.374274563e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.074599858e-07 wvoff=2.487297736e-08 pvoff=-1.983902501e-13 nfactor=-5.988435527e-01 lnfactor=2.807076281e-05 wnfactor=3.365484891e-06 pnfactor=-2.684356520e-11 eta0=0.08 etab=-0.07 u0=6.354263526e-02 lu0=-2.788507815e-07 wu0=-3.343222621e-08 pu0=2.666599830e-13 ua=2.585157423e-09 lua=-2.589886353e-14 wua=-3.105089609e-15 pua=2.476661701e-20 ub=-5.311598759e-19 lub=1.514413689e-23 wub=1.815674345e-24 pub=-1.448206551e-29 uc=-1.625786688e-10 luc=1.502525906e-15 wuc=1.801421739e-16 puc=-1.436838478e-21 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.373945912e+00 la0=-8.074969904e-08 wa0=-9.681314824e-09 pa0=7.721948369e-14 ags=3.469876285e-01 lags=-1.500014868e-08 wags=-1.798411182e-09 pags=1.434437218e-14 a1=0.0 a2=0.42385546 b0=-1.932656459e-07 lb0=1.541513076e-12 wb0=1.848164584e-13 pb0=-1.474121208e-18 b1=-3.240480314e-08 lb1=2.584651169e-13 wb1=3.098812995e-14 pb1=-2.471655389e-19 keta=2.343047201e-02 lketa=-1.991149009e-07 wketa=-2.387246100e-08 pketa=1.904099956e-13 dwg=0.0 dwb=0.0 pclm=6.357564328e-01 lpclm=-4.404625155e-06 wpclm=-5.280832413e-07 ppclm=4.212063752e-12 pdiblc1=0.39 pdiblc2=2.129425593e-02 lpdiblc2=-1.447180802e-07 wpdiblc2=-1.735066894e-08 ppdiblc2=1.383912952e-13 pdiblcb=-2.039148028e+01 lpdiblcb=1.449497539e-04 wpdiblcb=1.737844497e-05 ppdiblcb=-1.386128405e-10 drout=0.56 pscbe1=5.206373459e+09 lpscbe1=-3.545280514e+04 wpscbe1=-4.250539284e+03 ppscbe1=3.390287940e-2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.430167130e-01 lkt1=4.030876957e-07 wkt1=4.832734896e-08 pkt1=-3.854655078e-13 kt2=5.294212413e-02 lkt2=-5.868743411e-07 wkt2=-7.036206111e-08 pkt2=5.612173686e-13 at=-1.499647466e+05 lat=2.312798254e+00 wat=2.772880678e-01 pat=-2.211687340e-6 ute=-2.715155024e+00 lute=1.138557540e-05 wute=1.365049545e-06 pute=-1.088782082e-11 ua1=3.280622859e-09 lua1=-1.537019640e-14 wua1=-1.842777273e-15 pua1=1.469824215e-20 ub1=-4.028858998e-18 lub1=2.462072861e-23 wub1=2.951850319e-24 pub1=-2.354435960e-29 uc1=-5.067993504e-10 luc1=3.847616440e-15 wuc1=4.613018565e-16 puc1=-3.679406344e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.65 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.223228346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.818707001e-8 k1=4.568785944e-01 lk1=1.327020504e-7 k2=9.340993149e-03 lk2=-6.786532205e-08 pk2=2.081668171e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.167922808e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.287101972e-8 nfactor=2.949426389e+00 lnfactor=-2.307208158e-7 eta0=0.08 etab=-0.07 u0=2.924273440e-02 lu0=-5.270107433e-9 ua=-6.247801648e-10 lua=-2.959647776e-16 ub=1.360332146e-18 lub=5.733927629e-26 uc=2.621848235e-11 luc=-3.345848257e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.492475844e+00 la0=-1.026160561e-6 ags=3.537531077e-01 lags=-6.896253114e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.275941100e-02 lketa=8.954052784e-08 wketa=-3.469446952e-24 pketa=-6.938893904e-30 dwg=0.0 dwb=0.0 pclm=-3.634155134e-01 lpclm=3.564906175e-06 wpclm=1.110223025e-22 pdiblc1=0.39 pdiblc2=2.957262709e-03 lpdiblc2=1.540271552e-9 pdiblcb=-4.399015674e+00 lpdiblcb=1.739168118e-5 drout=0.56 pscbe1=7.777019419e+08 lpscbe1=-1.291188214e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912573382e-01 lkt1=-9.752116958e-9 kt2=-2.057529825e-02 lkt2=-4.893818432e-10 at=140000.0 ute=-1.488693675e+00 lute=1.603152885e-6 ua1=1.252307935e-09 lua1=8.079192830e-16 ub1=-9.358870489e-19 lub1=-4.923629781e-26 uc1=-3.049530213e-11 luc1=4.855057335e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.66 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.093723706e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.967987643e-8 k1=4.416709045e-01 lk1=1.931698936e-7 k2=1.666314832e-02 lk2=-9.697920683e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.640889714e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.793744597e-8 nfactor=3.384272625e+00 lnfactor=-1.959728587e-06 wnfactor=3.552713679e-21 eta0=0.08 etab=-0.07 u0=2.924253632e-02 lu0=-5.269319858e-9 ua=-2.473648295e-10 lua=-1.796619479e-15 ub=8.224210119e-19 lub=2.196147102e-24 uc=-2.997348756e-12 luc=1.128202696e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.427763872e+00 la0=-7.688569563e-7 ags=1.771075391e-01 lags=6.334042736e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.814126858e-02 lketa=-7.308613666e-08 wketa=1.387778781e-23 dwg=0.0 dwb=0.0 pclm=5.095155328e-01 lpclm=9.401361739e-8 pdiblc1=0.39 pdiblc2=1.415661641e-03 lpdiblc2=7.669887058e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.911105335e+08 lpscbe1=2.151803947e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.957157780e-01 lkt1=7.975246273e-9 kt2=-2.366218282e-02 lkt2=1.178449104e-8 at=1.684563584e+05 lat=-1.131463511e-1 ute=-1.740618726e+00 lute=2.604841151e-6 ua1=-6.739841536e-10 lua1=8.467118605e-15 pua1=-3.308722450e-36 ub1=8.183264192e-19 lub1=-7.024227620e-24 pub1=-3.081487911e-45 uc1=-6.492586981e-12 luc1=-4.688748644e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.67 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.269636961e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.491702467e-8 k1=5.981414663e-01 lk1=-1.160372166e-7 k2=-5.041999168e-02 lk2=3.558620112e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.009647561e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.917308910e-8 nfactor=2.817502433e+00 lnfactor=-8.397136079e-7 eta0=1.556199869e-01 leta0=-1.494353785e-7 etab=-5.596804500e-02 letab=-2.772905143e-8 u0=2.859798223e-02 lu0=-3.995593312e-9 ua=-9.275965507e-10 lua=-4.523890865e-16 ub=1.780184404e-18 lub=3.034763837e-25 uc=3.842701720e-11 luc=3.096008872e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.023864000e+04 lvsat=1.928977490e-2 a0=1.415845595e+00 la0=-7.453048199e-7 ags=3.271776224e-01 lags=3.368453795e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.678710971e-02 lketa=3.545980911e-08 wketa=1.387778781e-23 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=4.290014341e-01 lpclm=2.531204263e-7 pdiblc1=4.400712671e-01 lpdiblc1=-9.894763339e-8 pdiblc2=4.799318577e-03 lpdiblc2=9.833207738e-10 pdiblcb=-1.209086295e-03 lpdiblcb=-4.701408105e-8 drout=7.188175127e-01 ldrout=-3.138450042e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.117136320e-08 lalpha0=-2.314772989e-15 alpha1=9.993488080e-01 lalpha1=-2.951335560e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.258838054e-01 lkt1=6.759137127e-8 kt2=3.871048534e-04 lkt2=-3.574017210e-8 at=1.360768260e+05 lat=-4.915999135e-02 wat=-1.164153218e-16 ute=1.869609889e-01 lute=-1.204318517e-6 ua1=5.918675958e-09 lua1=-4.560874379e-15 ub1=-4.657704193e-18 lub1=3.797153610e-24 uc1=-7.733386419e-11 luc1=9.310451173e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.68 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.870056768e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.692114131e-9 k1=3.990662161e-01 lk1=7.828730192e-8 k2=6.570711535e-03 lk2=-2.004447595e-08 pk2=-6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.091905561e-01 ldsub=4.959692731e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.569585476e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.484466620e-9 nfactor=8.436487450e-01 lnfactor=1.087036036e-6 eta0=-4.616714939e-01 leta0=4.531250584e-07 weta0=5.898059818e-23 peta0=-1.162264729e-28 etab=-1.644253650e-01 letab=7.814004309e-8 u0=2.685234983e-02 lu0=-2.291618679e-9 ua=-1.301021280e-09 lua=-8.787576494e-17 ub=2.214008792e-18 lub=-1.199952198e-25 uc=6.310099629e-11 luc=6.874929471e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=5.704996039e+04 lvsat=3.216371986e-2 a0=-1.549019290e-01 la0=7.879583848e-7 ags=2.695021758e-01 lags=3.931444592e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.875782245e-02 lketa=-3.828231879e-08 wketa=-1.387778781e-23 pketa=-6.938893904e-30 dwg=0.0 dwb=0.0 pclm=8.676323403e-01 lpclm=-1.750429920e-07 wpclm=8.881784197e-22 pdiblc1=5.259075539e-01 lpdiblc1=-1.827355231e-7 pdiblc2=9.807043116e-03 lpdiblc2=-3.904899426e-9 pdiblcb=-7.258182741e-02 lpdiblcb=2.265542098e-8 drout=-1.766347053e-01 ldrout=5.602381421e-07 pdrout=-2.220446049e-28 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.765727360e-08 lalpha0=1.115456377e-15 alpha1=5.513023840e-01 lalpha1=1.422206881e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.431915482e-01 lkt1=-1.312751794e-8 kt2=-3.610930687e-02 lkt2=-1.147107452e-10 at=1.196012296e+05 lat=-3.307756865e-2 ute=-8.762049469e-01 lute=-1.665239728e-7 ua1=1.391698507e-09 lua1=-1.419287174e-16 ub1=-8.515011762e-19 lub1=8.178182225e-26 uc1=-2.098513587e-12 luc1=1.966457754e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.69 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.210479312e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.990085699e-8 k1=2.527004922e-01 lk1=1.479772922e-7 k2=5.872651086e-02 lk2=-4.487772962e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.819493130e-01 ldsub=6.256746383e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413312e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.155535806e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.422992879e-8 nfactor=3.861524120e+00 lnfactor=-3.498830736e-07 wnfactor=-3.552713679e-21 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.920295691e-02 letab=-1.881473159e-08 wetab=1.387778781e-23 petab=5.854691731e-30 u0=1.936882429e-02 lu0=1.271557234e-9 ua=-1.768133457e-09 lua=1.345331586e-16 ub=2.117932481e-18 lub=-7.424982916e-26 uc=6.395374912e-11 luc=6.468903149e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.097462453e+04 lvsat=1.601096598e-2 a0=1.5 ags=9.551765888e-01 lags=6.667018692e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=1.494316756e-02 lketa=-2.218194427e-8 dwg=0.0 dwb=0.0 pclm=7.364749379e-01 lpclm=-1.125942310e-7 pdiblc1=-5.222503249e-02 lpdiblc1=9.253421406e-8 pdiblc2=-4.545350845e-03 lpdiblc2=2.928792025e-09 ppdiblc2=4.336808690e-31 pdiblcb=4.582196898e-02 lpdiblcb=-3.372088902e-08 ppdiblcb=-6.938893904e-30 drout=1.449262890e+00 ldrout=-2.139102352e-7 pscbe1=8.077610961e+08 lpscbe1=-3.695337236e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.759816960e-08 lalpha0=-3.617762081e-15 alpha1=0.85 beta0=1.344390976e+01 lbeta0=1.981155425e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.977194842e-01 lkt1=1.283519537e-8 kt2=-4.310833573e-02 lkt2=3.217778860e-9 at=6.949658549e+04 lat=-9.220943808e-3 ute=-1.141734153e+00 lute=-4.009595862e-8 ua1=2.104407137e-09 lua1=-4.812749535e-16 ub1=-1.934788051e-18 lub1=5.975737015e-25 wub1=-7.703719778e-40 pub1=1.925929944e-46 uc1=-5.847484063e-11 luc1=4.650737639e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.70 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.170607816e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.899921892e-8 k1=0.90707349 k2=-1.569578983e-01 lk2=3.896279940e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586410187e-01 ldsub=-2.491733918e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-1.136835600e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280776e-8 nfactor=4.637117428e+00 lnfactor=-5.252726419e-7 eta0=6.941427212e-04 leta0=-6.153674857e-16 etab=-0.043998 u0=2.216395399e-02 lu0=6.394777856e-10 ua=-1.162846800e-09 lua=-2.343944841e-18 ub=1.468666835e-18 lub=7.257250696e-26 uc=5.323603314e-11 luc=8.892564569e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.251510632e+05 lvsat=8.282442839e-3 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.816207447e-01 lketa=2.226823259e-8 dwg=0.0 dwb=0.0 pclm=4.814953109e-01 lpclm=-5.493415810e-08 wpclm=-4.440892099e-22 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.16e-8 alpha1=0.85 beta0=1.485532343e+01 lbeta0=-1.210558988e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.24096074 kt2=-0.028878939 at=-4.265597014e+04 lat=1.614078651e-2 ute=-1.3190432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.71 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=8.4e-07 wmax=1.0e-6 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.112311471e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.313819688e-08 wvth0=1.700483939e-07 pvth0=-2.655067602e-14 k1=0.90707349 k2=-9.208700750e-02 lk2=-6.232401474e-09 wk2=-5.245945226e-08 pk2=8.190809038e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587284293e-01 ldsub=-1.613967235e-11 wdsub=-9.885022130e-11 pdsub=1.543407815e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-1.665995528e+01 lnfactor=2.799967102e-06 wnfactor=1.073285287e-05 pnfactor=-1.675784716e-12 eta0=-1.383068870e-02 leta0=2.267848679e-09 weta0=1.388983239e-08 peta0=-2.168702870e-15 etab=-0.043998 u0=2.657082505e-02 lu0=-4.859343515e-11 wu0=-4.122094249e-10 pu0=6.436073076e-17 ua=-1.268375502e-09 lua=1.413288451e-17 wua=8.584361323e-17 pua=-1.340327840e-23 ub=8.366006974e-18 lub=-1.004350593e-24 wub=-5.776708883e-24 pub=9.019522181e-31 uc=1.487513236e-10 luc=-6.020810825e-18 wuc=8.040084801e-17 puc=-1.255346681e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.553423676e+05 lvsat=-1.204510666e-02 wvsat=-8.495316084e-02 pvsat=1.326424672e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-7.679508232e-01 lketa=1.138154657e-07 wketa=5.402744889e-07 pketa=-8.435629760e-14 dwg=0.0 dwb=0.0 pclm=9.659855716e-02 lpclm=5.162081439e-09 wpclm=3.161606268e-08 ppclm=-4.936405563e-15 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.371808000e-08 lalpha0=5.514423739e-15 alpha1=0.85 beta0=1.923203543e+01 lbeta0=-8.044182041e-07 wbeta0=-4.002033251e-06 pbeta0=6.248614637e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-7.435506831e-01 lkt1=7.847238336e-08 wkt1=4.002033251e-07 pkt1=-6.248614637e-14 kt2=-0.028878939 at=4.168356834e+05 lat=-5.560240230e-02 wat=-2.601321613e-01 pat=4.061599514e-8 ute=-2.727950088e-01 lute=-1.633570076e-07 wute=-1.000508313e-06 pute=1.562153659e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.72 nmos lmin=2.0e-05 lmax=0.0001 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.73 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.634895033e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.074497225e-7 k1=6.308143008e-01 lk1=-1.254632799e-6 k2=-6.127234930e-02 lk2=4.953563007e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.061910635e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.168573159e-8 nfactor=3.627655214e+00 lnfactor=-5.640366163e-6 eta0=0.08 etab=-0.07 u0=2.155722531e-02 lu0=5.603055831e-8 ua=-1.314327444e-09 lua=5.203958101e-15 ub=1.749030239e-18 lub=-3.042969578e-24 uc=6.365044836e-11 luc=-3.019082999e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.361787763e+00 la0=1.622534711e-8 ags=3.447291181e-01 lags=3.014037474e-9 a1=0.0 a2=0.42385546 b0=3.883360838e-08 lb0=-3.097421418e-13 b1=6.511221529e-09 lb1=-5.193438844e-14 keta=-6.549435865e-03 lketa=4.000892163e-8 dwg=0.0 dwb=0.0 pclm=-2.742977677e-02 lpclm=8.850382462e-07 ppclm=-2.220446049e-28 pdiblc1=0.39 pdiblc2=-4.953474300e-04 lpdiblc2=2.907875958e-08 ppdiblc2=1.387778781e-29 pdiblcb=1.433005225e+00 lpdiblcb=-2.912531065e-05 wpdiblcb=5.551115123e-23 ppdiblcb=-6.439293543e-27 drout=0.56 pscbe1=-1.316089196e+08 lpscbe1=7.123668276e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.823254642e-01 lkt1=-8.099395856e-8 kt2=-3.542112043e-02 lkt2=1.179229150e-7 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.000875981e+00 lute=-2.287747387e-6 ua1=9.663958972e-10 lua1=3.088392584e-15 ub1=-3.218176240e-19 lub1=-4.947137544e-24 uc1=7.252035853e-11 luc1=-7.731163462e-16 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.74 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.223228346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.818707001e-8 k1=4.568785944e-01 lk1=1.327020504e-7 k2=9.340993149e-03 lk2=-6.786532205e-08 wk2=1.734723476e-24 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.167922808e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=4.287101972e-8 nfactor=2.949426389e+00 lnfactor=-2.307208158e-7 eta0=0.08 etab=-0.07 u0=2.924273440e-02 lu0=-5.270107433e-9 ua=-6.247801648e-10 lua=-2.959647776e-16 ub=1.360332146e-18 lub=5.733927629e-26 uc=2.621848235e-11 luc=-3.345848257e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.492475844e+00 la0=-1.026160561e-6 ags=3.537531077e-01 lags=-6.896253114e-8 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.275941100e-02 lketa=8.954052784e-08 wketa=3.469446952e-24 pketa=-1.387778781e-29 dwg=0.0 dwb=0.0 pclm=-3.634155134e-01 lpclm=3.564906175e-06 wpclm=2.220446049e-22 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=2.957262709e-03 lpdiblc2=1.540271552e-9 pdiblcb=-4.399015674e+00 lpdiblcb=1.739168118e-5 drout=0.56 pscbe1=7.777019419e+08 lpscbe1=-1.291188214e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.912573382e-01 lkt1=-9.752116958e-9 kt2=-2.057529825e-02 lkt2=-4.893818432e-10 at=140000.0 ute=-1.488693675e+00 lute=1.603152885e-6 ua1=1.252307935e-09 lua1=8.079192830e-16 ub1=-9.358870489e-19 lub1=-4.923629781e-26 uc1=-3.049530213e-11 luc1=4.855057335e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.75 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.093723706e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.967987643e-8 k1=4.416709045e-01 lk1=1.931698936e-7 k2=1.666314832e-02 lk2=-9.697920683e-08 pk2=2.775557562e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.640889714e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-7.793744597e-8 nfactor=3.384272625e+00 lnfactor=-1.959728587e-6 eta0=0.08 etab=-0.07 u0=2.924253632e-02 lu0=-5.269319858e-9 ua=-2.473648295e-10 lua=-1.796619479e-15 ub=8.224210119e-19 lub=2.196147102e-24 uc=-2.997348756e-12 luc=1.128202696e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.427763872e+00 la0=-7.688569563e-7 ags=1.771075391e-01 lags=6.334042736e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.814126858e-02 lketa=-7.308613666e-08 wketa=-1.387778781e-23 pketa=-2.775557562e-29 dwg=0.0 dwb=0.0 pclm=5.095155328e-01 lpclm=9.401361739e-8 pdiblc1=0.39 pdiblc2=1.415661641e-03 lpdiblc2=7.669887058e-9 pdiblcb=-0.025 drout=0.56 pscbe1=6.911105335e+08 lpscbe1=2.151803947e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.957157780e-01 lkt1=7.975246273e-9 kt2=-2.366218282e-02 lkt2=1.178449104e-8 at=1.684563584e+05 lat=-1.131463511e-1 ute=-1.740618726e+00 lute=2.604841151e-6 ua1=-6.739841536e-10 lua1=8.467118605e-15 ub1=8.183264192e-19 lub1=-7.024227620e-24 pub1=3.081487911e-45 uc1=-6.492586981e-12 luc1=-4.688748644e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.76 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.269636961e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.491702467e-8 k1=5.981414663e-01 lk1=-1.160372166e-7 k2=-5.041999168e-02 lk2=3.558620112e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.009647561e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-4.917308910e-8 nfactor=2.817502433e+00 lnfactor=-8.397136079e-7 eta0=1.556199869e-01 leta0=-1.494353785e-7 etab=-5.596804500e-02 letab=-2.772905143e-8 u0=2.859798223e-02 lu0=-3.995593312e-9 ua=-9.275965507e-10 lua=-4.523890865e-16 ub=1.780184404e-18 lub=3.034763837e-25 uc=3.842701720e-11 luc=3.096008872e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.023864000e+04 lvsat=1.928977490e-2 a0=1.415845595e+00 la0=-7.453048199e-7 ags=3.271776224e-01 lags=3.368453795e-7 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.678710971e-02 lketa=3.545980911e-8 dwg=0.0 dwb=0.0 pclm=4.290014341e-01 lpclm=2.531204263e-7 pdiblc1=4.400712671e-01 lpdiblc1=-9.894763339e-8 pdiblc2=4.799318577e-03 lpdiblc2=9.833207738e-10 pdiblcb=-1.209086295e-03 lpdiblcb=-4.701408105e-8 drout=7.188175127e-01 ldrout=-3.138450042e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.117136320e-08 lalpha0=-2.314772989e-15 alpha1=9.993488080e-01 lalpha1=-2.951335560e-7 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.258838054e-01 lkt1=6.759137127e-8 kt2=3.871048534e-04 lkt2=-3.574017210e-8 at=1.360768260e+05 lat=-4.915999135e-2 ute=1.869609889e-01 lute=-1.204318517e-6 ua1=5.918675958e-09 lua1=-4.560874379e-15 ub1=-4.657704193e-18 lub1=3.797153610e-24 uc1=-7.733386419e-11 luc1=9.310451173e-17 puc1=-5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.77 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.955018131e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.562810135e-08 wvth0=7.286287958e-08 pvth0=-7.112407982e-14 k1=-1.877614812e-01 lk1=6.511109430e-07 wk1=4.672803325e-07 pk1=-4.561291546e-13 k2=1.683158353e-01 lk2=-1.779297141e-07 wk2=-1.287947306e-07 pk2=1.257211732e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.889748954e-01 ldsub=6.933016149e-08 wdsub=1.609736674e-08 pdsub=-1.571321918e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.450009742e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.187751262e-09 wvoff=-9.521600473e-09 pvoff=9.294376999e-15 nfactor=-1.073338238e-01 lnfactor=2.015324357e-06 wnfactor=7.572503019e-07 pnfactor=-7.391792807e-13 eta0=-4.616714938e-01 leta0=4.531250583e-07 weta0=-1.059644698e-16 peta0=1.034357981e-22 etab=-1.664973958e-01 letab=8.016262691e-08 wetab=1.649920800e-09 petab=-1.610547090e-15 u0=3.316325832e-02 lu0=-8.451923647e-09 wu0=-5.025262832e-09 pu0=4.905339960e-15 ua=-1.077074867e-09 lua=-3.064779208e-16 wua=-1.783244976e-16 pua=1.740689618e-22 ub=1.779380939e-18 lub=3.042606742e-25 wub=3.460863361e-25 pub=-3.378273318e-31 uc=-1.026813584e-10 luc=1.687010541e-16 wuc=1.320095050e-16 puc=-1.288592301e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=4.676203749e+05 lvsat=-3.686088423e-01 wvsat=-3.269298308e-01 pvsat=3.191279773e-7 a0=-9.200614575e-01 la0=1.534858146e-06 wa0=6.092827597e-07 pa0=-5.947428360e-13 ags=-5.956204410e+00 lags=6.470280783e-06 wags=4.957418091e-06 pags=-4.839114266e-12 a1=0.0 a2=0.42385546 b0=1.213199662e-16 lb0=-1.184247865e-22 wb0=-9.660490534e-23 pb0=9.429952588e-29 b1=-9.314584709e-18 lb1=9.092301459e-24 wb1=7.417036141e-24 pb1=-7.240035991e-30 keta=2.114101305e-01 lketa=-1.970530922e-07 wketa=-1.295171052e-07 pketa=1.264263090e-13 dwg=0.0 dwb=0.0 pclm=5.481086146e-01 lpclm=1.368556195e-07 wpclm=2.544309914e-07 ppclm=-2.483592502e-13 pdiblc1=-1.973953426e-01 lpdiblc1=5.233064731e-07 wpdiblc1=5.759530771e-07 ppdiblc1=-5.622085328e-13 pdiblc2=-5.324133019e-04 lpdiblc2=6.187816203e-09 wpdiblc2=8.233123035e-09 ppdiblc2=-8.036647787e-15 pdiblcb=-5.340990697e-01 lpdiblcb=4.731590158e-07 wpdiblcb=3.674978727e-07 ppdiblcb=-3.587279035e-13 drout=-1.766353686e-01 ldrout=5.602387895e-07 wdrout=5.281445228e-13 pdrout=-5.155408820e-19 pscbe1=-1.607222313e+09 lpscbe1=2.349776360e+03 wpscbe1=1.916827798e+03 ppscbe1=-1.871084619e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.568768658e-05 lalpha0=-2.504656291e-11 walpha0=-2.043261945e-11 palpha0=1.994501542e-17 alpha1=5.513023840e-01 lalpha1=1.422206881e-7 beta0=4.142961286e+01 lbeta0=-2.691169162e-05 wbeta0=-2.195318647e-05 pbeta0=2.142929563e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.974760364e-01 lkt1=3.986152520e-08 wkt1=4.322576081e-08 pkt1=-4.219422125e-14 kt2=-3.855180350e-02 lkt2=2.269498146e-09 wkt2=1.944916102e-09 pkt2=-1.898502624e-15 at=-1.421385482e+05 lat=2.224160511e-01 wat=2.084186737e-01 pat=-2.034449705e-7 ute=-1.435378758e+00 lute=3.793057145e-07 wute=4.452600407e-07 pute=-4.346343550e-13 ua1=-3.451243119e-10 lua1=1.553446562e-15 wua1=1.383000748e-15 pua1=-1.349996818e-21 ub1=-5.341608751e-19 lub1=-2.279854699e-25 wub1=-2.526923696e-25 pub1=2.466621189e-31 uc1=-2.239642498e-10 luc1=2.362357099e-16 wuc1=1.766676922e-16 puc1=-1.724516944e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.78 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='7.019307173e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.266013141e-08 wvth0=-6.440550672e-08 pvth0=-5.765659441e-15 k1=1.426355886e+00 lk1=-1.174284437e-07 wk1=-9.345606642e-07 pk1=2.113378102e-13 k2=-2.731314950e-01 lk2=3.225925199e-08 wk2=2.642525566e-07 pk2=-6.142278999e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.223806346e-01 ldsub=5.342448646e-08 wdsub=-3.219473359e-08 pdsub=7.280388301e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413304e-03 lcdscd=-1.441936597e-09 wcdscd=6.155763399e-18 pcdscd=-2.930981846e-24 cit=0.0 voff='-1.394687272e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.821853256e-09 wvoff=1.904320076e-08 pvoff=-4.306353200e-15 nfactor=5.763489260e+00 lnfactor=-7.799858629e-07 wnfactor=-1.514500605e-06 pnfactor=3.424831092e-13 eta0=9.325986799e-01 leta0=-2.107371651e-07 weta0=-5.891998001e-17 peta0=8.103628879e-23 etab=4.334701840e-02 letab=-1.975185307e-08 wetab=-3.299841571e-09 petab=7.462129661e-16 u0=1.667671323e-02 lu0=-6.020860148e-10 wu0=2.143679585e-09 pu0=1.491948394e-15 ua=-2.216026280e-09 lua=2.358178492e-16 wua=3.566489928e-16 pua=-8.065117599e-23 ub=2.987188189e-18 lub=-2.708198382e-25 wub=-6.921726734e-25 pub=1.565251600e-31 uc=3.955184586e-10 luc=-6.850981403e-17 wuc=-2.640190100e-16 puc=5.970420287e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.277956344e+05 lvsat=1.529581547e-01 wvsat=5.723438193e-01 pvsat=-1.090485814e-7 a0=3.030319055e+00 la0=-3.460602291e-07 wa0=-1.218565517e-06 pa0=2.755615313e-13 ags=1.340658976e+01 lags=-2.749042582e-06 wags=-9.914836182e-06 pags=2.242101395e-12 a1=0.0 a2=0.42385546 b0=-2.426399324e-16 lb0=5.486962376e-23 wb0=1.932098107e-22 pb0=-4.369169375e-29 b1=1.862916942e-17 lb1=-4.212725855e-24 wb1=-1.483407228e-23 pb1=3.354517770e-30 keta=-3.103614485e-01 lketa=5.138114037e-08 wketa=2.590342103e-07 pketa=-5.857696016e-14 dwg=0.0 dwb=0.0 pclm=1.375522390e+00 lpclm=-2.571058657e-07 wpclm=-5.088619830e-07 ppclm=1.150720135e-13 pdiblc1=1.394380761e+00 lpdiblc1=-2.345954338e-07 wpdiblc1=-1.151906154e-06 ppdiblc1=2.604874502e-13 pdiblc2=1.613356198e-02 lpdiblc2=-1.747454603e-09 wpdiblc2=-1.646624606e-08 ppdiblc2=3.723611017e-15 pdiblcb=9.688564536e-01 lpdiblcb=-2.424522152e-07 wpdiblcb=-7.349957455e-07 ppdiblcb=1.662089979e-13 drout=1.449264214e+00 ldrout=-2.139105341e-07 wdrout=-1.054410701e-12 pdrout=2.379706321e-19 pscbe1=5.622205722e+09 lpscbe1=-1.092414587e+03 wpscbe1=-3.833655595e+03 ppscbe1=8.669275417e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.128246043e-05 lalpha0=1.160169501e-11 walpha0=4.086523891e-11 palpha0=-9.241101665e-18 alpha1=0.85 beta0=-4.169531597e+01 lbeta0=1.266707949e-05 wbeta0=4.390637294e-05 pbeta0=-9.928811551e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.891505079e-01 lkt1=-1.171615863e-08 wkt1=-8.645152155e-08 pkt1=1.954980126e-14 kt2=-3.822334249e-02 lkt2=2.113106030e-09 wkt2=-3.889832193e-09 pkt2=8.796310899e-16 at=5.929761411e+05 lat=-1.275985166e-01 wat=-4.168373475e-01 pat=9.426193042e-8 ute=-2.338653081e-02 lute=-2.929946166e-07 wute=-8.905200814e-07 pute=2.013786492e-13 ua1=5.578052773e-09 lua1=-1.266791282e-15 wua1=-2.766001494e-15 pua1=6.254925134e-22 ub1=-2.569468657e-18 lub1=7.410978359e-25 wub1=5.053847423e-25 pub1=-1.142856848e-31 uc1=3.852566319e-10 luc1=-5.383628390e-17 wuc1=-3.533353844e-16 puc1=7.990185051e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.79 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='8.841191988e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.385950585e-08 wvth0=-2.126538106e-07 pvth0=2.775861900e-14 k1=9.070734930e-01 lk1=-4.748850202e-16 wk1=-2.421877809e-15 pk1=3.781419622e-22 k2=-1.581819230e-01 lk2=6.265015584e-09 wk2=9.746688340e-10 pk2=-1.886181556e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.587177398e-01 ldsub=-1.984115670e-11 wdsub=-6.109158814e-11 pdsub=1.381503307e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000031e-03 lcdscd=-5.025100128e-18 wcdscd=-2.450002701e-17 pcdscd=4.001398171e-24 cit=0.0 voff='-1.136835613e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280753e-08 wvoff=9.995093642e-16 pvoff=-1.791236048e-22 nfactor=2.330204247e+01 lnfactor=-4.746084131e-06 wnfactor=-1.486254384e-05 pnfactor=3.360956214e-12 eta0=-1.008629497e-02 leta0=2.437844358e-09 weta0=8.584268489e-09 peta0=-1.941212071e-15 etab=-4.399799987e-02 letab=-2.050434822e-17 wetab=-1.045705744e-16 petab=1.632724511e-23 u0=3.008992169e-02 lu0=-3.635295323e-09 wu0=-6.311305412e-09 pu0=3.403924881e-15 ua=-1.214258677e-09 lua=9.282130514e-18 wua=4.093835200e-17 pua=-9.257634536e-24 ub=2.675122220e-18 lub=-2.002504882e-25 wub=-9.606787065e-25 pub=2.172440403e-31 uc=-4.621647650e-10 luc=1.254432394e-16 wuc=4.104043783e-16 puc=-9.280720448e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.181362131e+05 lvsat=3.770581185e-02 wvsat=1.937252790e-01 pvsat=-2.342929912e-8 a0=1.500000009e+00 la0=-1.450684017e-15 wa0=-7.398387680e-15 pa0=1.155153306e-21 ags=1.250000002e+00 lags=-3.106048752e-16 wags=-1.584059106e-15 pags=2.473292682e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=4.747288614e-03 lketa=-1.987628900e-08 wketa=-1.484015103e-07 pketa=3.355892394e-14 dwg=0.0 dwb=0.0 pclm=1.253453660e+00 lpclm=-2.295017314e-07 wpclm=-6.146965380e-07 ppclm=1.390050164e-13 pdiblc1=3.569721484e-01 lpdiblc1=2.483540040e-16 wpdiblc1=1.266587724e-15 ppdiblc1=-1.977599196e-22 pdiblc2=8.406112143e-03 lpdiblc2=-6.658944229e-18 wpdiblc2=-3.396011250e-17 ppdiblc2=5.302397410e-24 pdiblcb=-1.032957699e-01 lpdiblcb=-1.971667274e-17 wpdiblcb=-1.005533434e-16 ppdiblcb=1.569999686e-23 drout=5.033266684e-01 ldrout=-1.315386911e-15 wdrout=-6.708376077e-15 pdrout=1.047419040e-21 pscbe1=7.914198808e+08 lpscbe1=-1.299495697e-07 wpscbe1=-6.627311707e-07 ppscbe1=1.034765244e-13 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.520576188e-07 lalpha0=-2.950116442e-14 walpha0=-1.038810536e-13 palpha0=2.349124621e-20 alpha1=0.85 beta0=1.148724706e+01 lbeta0=6.405874201e-07 wbeta0=2.681938591e-06 pbeta0=-6.064828653e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-9.585292216e-02 lkt1=-3.281410148e-08 wkt1=-1.155467434e-07 pkt1=2.612927835e-14 kt2=-2.887893895e-02 lkt2=-7.882083874e-18 wkt2=-4.019806710e-17 pkt2=6.276368314e-24 at=-1.513706568e+05 lat=4.072509088e-02 wat=8.656754808e-02 pat=-1.957603905e-8 ute=-1.268048809e+00 lute=-1.153166767e-08 wute=-4.060591577e-08 pute=9.182459393e-15 ua1=-2.384732647e-11 lua1=-1.487216600e-24 wua1=-7.584694177e-24 pua1=1.184243813e-30 ub1=7.077531835e-19 lub1=-2.112662719e-33 wub1=-1.077442402e-32 pub1=1.682275540e-39 uc1=1.471862498e-10 luc1=3.058996623e-26 wuc1=1.560062635e-25 puc1=-2.435824599e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.80 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=7.4e-07 wmax=8.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='8.450674508e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.776212212e-08 wvth0=-1.754076457e-07 pvth0=2.194315179e-14 k1=0.90707349 k2=-1.448299398e-01 lk2=4.180290326e-09 wk2=-1.046120466e-08 pk2=-1.006300131e-16 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.584252728e-01 ldsub=2.582347576e-11 wdsub=1.425478955e-10 pdsub=-1.798042135e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999993e-03 lcdscd=8.702153581e-19 wcdscd=5.565652106e-18 pcdscd=-6.929378946e-25 cit=0.0 voff='-2.075299990e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.217839163e-16 wvoff=-7.688072401e-16 pvoff=9.697420644e-23 nfactor=-4.482171118e+01 lnfactor=5.890486268e-06 wnfactor=3.315755219e-05 pnfactor=-4.136709499e-12 eta0=2.876702308e-02 leta0=-3.628556861e-09 weta0=-2.002995755e-08 peta0=2.526498726e-15 etab=-0.043998 u0=-6.292865836e-02 lu0=1.088825369e-08 wu0=7.085461823e-08 pu0=-8.644453773e-15 ua=-1.029853534e-09 lua=-1.951015083e-17 wua=-1.040871361e-16 pua=1.338606508e-23 ub=-3.284610577e-18 lub=7.302783517e-25 wub=3.500468162e-24 pub=-4.793015873e-31 uc=1.452323505e-09 luc=-1.734773010e-16 wuc=-9.576102154e-16 puc=1.207891221e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-2.889479130e+05 lvsat=6.437566743e-02 wvsat=3.484553924e-01 pvsat=-4.758824011e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.243131449e-01 lketa=6.272909085e-08 wketa=3.462701911e-07 pketa=-4.367713683e-14 dwg=0.0 dwb=0.0 pclm=-9.768628110e-01 lpclm=1.187309611e-07 wpclm=8.863940278e-07 ppclm=-9.536926020e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.181192019e-07 lalpha0=4.391036365e-14 walpha0=2.423891341e-13 palpha0=-3.057399582e-20 alpha1=0.85 beta0=1.955789333e+01 lbeta0=-6.195310072e-07 wbeta0=-4.261508034e-06 pbeta0=4.776391168e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.541912705e-01 lkt1=2.313541487e-08 wkt1=1.697916332e-07 pkt1=-1.842231442e-14 kt2=-0.028878939 at=3.438198224e+05 lat=-3.659196977e-02 wat=-2.019909455e-01 pat=2.547832990e-8 ute=-2.275028667e+00 lute=1.456941394e-07 wute=5.938343087e-07 pute=-8.987649950e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.81 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.82 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.292369027e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.191684330e-06 wvth0=2.384946925e-08 pvth0=-4.764202412e-13 k1=7.553195353e-01 lk1=-3.741766297e-06 wk1=-8.669075371e-08 pk1=1.731746286e-12 k2=-1.261738584e-01 lk2=1.791837673e-06 wk2=4.518975254e-08 pk2=-9.027166426e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.365377804e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.645244138e-07 wvoff=2.112987279e-08 pvoff=-4.220932124e-13 nfactor=3.370194296e+00 lnfactor=-4.972918408e-07 wnfactor=1.792654032e-07 pnfactor=-3.581030075e-12 eta0=0.08 etab=-0.07 u0=1.647114083e-02 lu0=1.576308735e-07 wu0=3.541349070e-09 pu0=-7.074247065e-14 ua=-1.802840015e-09 lua=1.496255165e-14 wua=3.401425097e-16 pua=-6.794733032e-21 ub=2.179925653e-18 lub=-1.165059497e-23 wub=-3.000247207e-25 pub=5.993334623e-30 uc=6.597431300e-11 luc=-3.483301360e-16 wuc=-1.618065118e-18 puc=3.232268885e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.165571201e+00 la0=3.935874094e-06 wa0=1.366220609e-07 pa0=-2.729180869e-12 ags=5.054877156e-01 lags=-3.208321569e-06 wags=-1.119333178e-07 pags=2.235995179e-12 a1=0.0 a2=0.42385546 b0=1.372239775e-07 lb0=-2.275201536e-12 wb0=-6.850744297e-14 pb0=1.368513998e-18 b1=1.531817597e-08 lb1=-2.278633082e-13 wb1=-6.132123855e-15 pb1=1.224961401e-19 keta=-3.274795282e-02 lketa=5.633540592e-07 wketa=1.824155578e-08 pketa=-3.643957991e-13 dwg=0.0 dwb=0.0 pclm=-1.467841810e-01 lpclm=3.269278057e-06 wpclm=8.310432329e-08 ppclm=-1.660103264e-12 pdiblc1=0.39 pdiblc2=-7.548456606e-03 lpdiblc2=1.699726277e-07 wpdiblc2=4.910952963e-09 ppdiblc2=-9.810186428e-14 pdiblcb=1.125480882e+01 lpdiblcb=-2.253269950e-04 wpdiblcb=-6.838745051e-06 ppdiblcb=1.366117012e-10 drout=0.56 pscbe1=-5.189850205e+08 lpscbe1=1.486194595e+04 wpscbe1=2.697230063e+02 ppscbe1=-5.388023456e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.763255054e-01 lkt1=-2.008499515e-07 wkt1=-4.177663310e-09 pkt1=8.345357045e-14 kt2=-3.512857767e-02 lkt2=1.120790409e-07 wkt2=-2.036922630e-10 pkt2=4.068984347e-15 at=1.982637300e+05 lat=-4.647194343e-1 ute=-8.996826457e-01 lute=-4.309199207e-06 wute=-7.045909762e-08 pute=1.407500517e-12 ua1=5.387868935e-10 lua1=1.163036820e-14 wua1=2.977364523e-16 pua1=-5.947623864e-21 ub1=8.810493406e-20 lub1=-1.313580631e-23 wub1=-2.854216986e-25 pub1=5.701622668e-30 uc1=9.414572346e-11 luc1=-1.205107577e-15 wuc1=-1.505735234e-17 puc1=3.007877181e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.83 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.921751317e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.079331442e-07 wvth0=-4.863689711e-08 pvth0=1.017408750e-13 k1=5.911392919e-01 lk1=-2.432242347e-06 wk1=-9.348330698e-08 pk1=1.785924615e-12 k2=-2.735954208e-02 lk2=1.003681247e-06 wk2=2.555392207e-08 pk2=-7.460985882e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.086682430e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.422331929e-07 wvoff=-5.656621301e-09 pvoff=-2.084404926e-13 nfactor=3.715913743e+00 lnfactor=-3.254797166e-06 wnfactor=-5.336913473e-07 pnfactor=2.105609929e-12 eta0=0.08 etab=-0.07 u0=5.298182253e-02 lu0=-1.335832891e-07 wu0=-1.652909976e-08 pu0=8.934215879e-14 ua=1.746990347e-09 lua=-1.335137810e-14 wua=-1.651421116e-15 pua=9.090249297e-21 ub=-4.422287084e-19 lub=9.264064832e-24 wub=1.255090677e-24 pub=-6.410477284e-30 uc=1.381727663e-10 luc=-9.241948184e-16 wuc=-7.795175273e-17 puc=6.411705627e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.051688700e+00 la0=-3.131919594e-06 wa0=-3.893698455e-07 pa0=1.466202111e-12 ags=3.051349040e-01 lags=-1.610280296e-06 wags=3.385198015e-08 pags=1.073191816e-12 a1=0.0 a2=0.42385546 b0=-7.292167675e-08 lb0=-5.990512180e-13 wb0=5.077405093e-14 pb0=4.171085802e-19 b1=-4.030522242e-09 lb1=-7.353545979e-14 wb1=2.806380088e-15 pb1=5.120141701e-20 keta=1.893225442e-02 lketa=1.511456978e-07 wketa=-2.206633618e-08 pketa=-4.289457096e-14 dwg=0.0 dwb=0.0 pclm=1.867328499e+00 lpclm=-1.279555860e-05 wpclm=-1.553226902e-06 ppclm=1.139149713e-11 pdiblc1=0.39 pdiblc2=3.394918562e-02 lpdiblc2=-1.610182104e-07 wpdiblc2=-2.157911807e-08 ppdiblc2=1.131865449e-13 pdiblcb=-3.386442646e+01 lpdiblcb=1.345501618e-04 wpdiblcb=2.051623515e-05 ppdiblcb=-8.157534117e-11 drout=0.56 pscbe1=1.711985740e+09 lpscbe1=-2.932580246e+03 wpscbe1=-6.505249915e+02 ppscbe1=1.951999728e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.248595398e-01 lkt1=1.862641072e-07 wkt1=2.339660812e-08 pkt1=-1.364825686e-13 kt2=-9.319538423e-02 lkt2=5.752277871e-07 wkt2=5.056405871e-08 pkt2=-4.008615018e-13 at=140000.0 ute=-3.224607310e+00 lute=1.423471610e-05 wute=1.208685418e-06 pute=-8.795130101e-12 ua1=-5.233895304e-10 lua1=2.010243181e-14 wua1=1.236386183e-15 pua1=-1.343442177e-20 ub1=-3.190224405e-19 lub1=-9.888503004e-24 wub1=-4.295117233e-25 pub1=6.850904301e-30 uc1=2.437299205e-10 luc1=-2.398211476e-15 wuc1=-1.909380865e-16 puc1=1.703636373e-21 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.84 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='3.324039326e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.249524725e-07 wvth0=1.232199380e-07 pvth0=-5.815852738e-13 k1=-3.497273802e-01 lk1=1.308771499e-06 wk1=5.510363804e-07 pk1=-7.767733172e-13 k2=3.963939237e-01 lk2=-6.812201634e-07 wk2=-2.643997038e-07 pk2=4.067964617e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.436826144e+00 ldsub=7.939652317e-06 wdsub=1.390354101e-06 pdsub=-5.528236994e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='2.560079898e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.107769105e-06 wvoff=-2.384187149e-07 pvoff=7.170532471e-13 nfactor=9.065216592e+00 lnfactor=-2.452435280e-05 wnfactor=-3.955539027e-06 pnfactor=1.571134168e-11 eta0=-4.491589281e-01 leta0=2.104007864e-06 weta0=3.684438368e-07 peta0=-1.464982803e-12 etab=3.925980567e-01 letab=-1.839352787e-06 wetab=-3.220987001e-07 petab=1.280708237e-12 u0=2.347866857e-02 lu0=-1.627473659e-08 wu0=4.013277368e-09 pu0=7.662873572e-15 ua=2.838977358e-09 lua=-1.769326696e-14 wua=-2.148964511e-15 pua=1.106854950e-20 ub=-4.919382610e-18 lub=2.706583764e-23 wub=3.997914510e-24 pub=-1.731631787e-29 uc=-2.628408164e-10 luc=6.702897242e-16 wuc=1.809243293e-16 puc=-3.881559468e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.960688333e-01 la0=4.246277360e-06 wa0=8.576070848e-07 pa0=-3.491947752e-12 ags=-8.312115197e-01 lags=2.907987628e-06 wags=7.020744109e-07 pags=-1.583751447e-12 a1=0.0 a2=0.42385546 b0=-4.345130239e-09 lb0=-8.717208933e-13 wb0=3.025435973e-15 pb0=6.069635671e-19 b1=8.800153735e-09 lb1=-1.245519724e-13 wb1=-6.127388643e-15 pb1=8.672329648e-20 keta=2.142250194e-01 lketa=-6.253648954e-07 wketa=-1.295667662e-07 pketa=3.845417587e-13 dwg=0.0 dwb=0.0 pclm=-3.578301750e+00 lpclm=8.857007879e-06 wpclm=2.846273593e-06 ppclm=-6.101515171e-12 pdiblc1=0.39 pdiblc2=-5.715063365e-03 lpdiblc2=-3.307762063e-09 wpdiblc2=4.964995469e-09 ppdiblc2=7.643539485e-15 pdiblcb=5.820108933e-02 lpdiblcb=-3.308188465e-07 wpdiblcb=-5.793142088e-08 ppdiblcb=2.303432081e-13 drout=0.56 pscbe1=1.146799543e+09 lpscbe1=-6.853230616e+02 wpscbe1=-3.172880548e+02 ppscbe1=6.270043475e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-5.449986400e-01 lkt1=1.061567109e-06 wkt1=1.735711697e-07 pkt1=-7.335970491e-13 kt2=-8.362615554e-02 lkt2=5.371792324e-07 wkt2=4.175183485e-08 pkt2=-3.658229013e-13 at=1.562757189e+05 lat=-6.471447193e-02 wat=8.481160017e-03 pat=-3.372224567e-8 ute=-7.581647527e+00 lute=3.155890056e-05 wute=4.067003215e-06 pute=-2.016019040e-11 ua1=-1.963254543e-08 lua1=9.608303450e-14 wua1=1.320050496e-14 pua1=-6.100538515e-20 ub1=1.634205074e-17 lub1=-7.613519586e-23 wub1=-1.080888982e-23 pub1=4.812072319e-29 uc1=-1.069321342e-10 luc1=-1.003931456e-15 wuc1=6.993424884e-17 puc1=6.663724895e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.85 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='8.114216701e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.165172333e-08 wvth0=-1.980629670e-07 pvth0=5.331344099e-14 k1=6.424935211e-01 lk1=-6.519919438e-07 wk1=-3.088153742e-08 pk1=3.731756294e-13 k2=-5.325272419e-02 lk2=2.073427648e-07 wk2=1.972380662e-09 pk2=-1.195910037e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.846493088e+00 ldsub=-4.477041017e-06 wdsub=-2.780708202e-06 pdsub=2.714349382e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.444927014e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.890192907e-08 wvoff=1.695641248e-07 pvoff=-8.917632980e-14 nfactor=-2.448385145e+00 lnfactor=-1.771909917e-06 wnfactor=3.666542735e-06 pnfactor=6.490715103e-13 eta0=1.213937514e+00 leta0=-1.182496888e-06 weta0=-7.368874447e-07 peta0=7.193021338e-13 etab=-9.811641583e-01 letab=8.753881819e-07 wetab=6.441974002e-07 petab=-6.288242734e-13 u0=1.338629348e-02 lu0=3.669169144e-09 wu0=1.059162506e-08 pu0=-5.336836133e-15 ua=-9.031842606e-09 lua=5.765087721e-15 wua=5.642840652e-15 pua=-4.329117186e-21 ub=1.335822209e-17 lub=-9.053194994e-24 wub=-8.061579233e-24 pub=6.514881860e-30 uc=-1.187470309e-10 luc=3.855408074e-16 wuc=1.094374606e-16 puc=-2.468881719e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.694418099e+04 lvsat=1.048455140e-01 wvsat=3.014515251e-02 pvsat=-5.957092110e-8 a0=7.598366558e+00 la0=-1.038166966e-05 wa0=-4.304778061e-06 pa0=6.709627380e-12 ags=4.408247860e+00 lags=-7.445896674e-06 wags=-2.841575747e-06 pags=5.418983202e-12 a1=0.0 a2=0.42385546 b0=-1.294931649e-07 lb0=-6.244113568e-13 wb0=9.016375983e-14 pb0=4.347663883e-19 b1=-9.267407280e-08 lb1=7.597489968e-14 wb1=6.452728876e-14 pb1=-5.289995510e-20 keta=-6.862209452e-01 lketa=1.154038791e-06 wketa=4.591519098e-07 pketa=-7.788464108e-13 dwg=0.0 dwb=0.0 pclm=2.310888861e+00 lpclm=-2.780833698e-06 wpclm=-1.310324341e-06 ppclm=2.112487645e-12 pdiblc1=5.430714416e-01 lpdiblc1=-3.024899864e-07 wpdiblc1=-7.171716755e-08 ppdiblc1=1.417228766e-13 pdiblc2=-2.758207008e-02 lpdiblc2=3.990441711e-08 wpdiblc2=2.254657805e-08 ppdiblc2=-2.710005880e-14 pdiblcb=1.557888629e-01 lpdiblcb=-5.236655591e-07 wpdiblcb=-1.093148461e-07 ppdiblcb=3.318838444e-13 drout=4.153991572e+00 ldrout=-7.102216130e-06 wdrout=-2.391849865e-06 pdrout=4.726620624e-12 pscbe1=3.653269851e+08 lpscbe1=8.589729929e+02 wpscbe1=3.026549961e+02 ppscbe1=-5.980874334e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.613969708e-05 lalpha0=-7.135767235e-11 walpha0=-2.514171650e-11 palpha0=4.968345108e-17 alpha1=2.005432075e+00 lalpha1=-2.283290919e-06 walpha1=-7.005176692e-07 palpha1=1.384318185e-12 beta0=3.755885028e+01 lbeta0=-4.683215121e-05 wbeta0=-1.650108287e-05 pbeta0=3.260838391e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=1.166165634e-01 lkt1=-2.458745130e-07 wkt1=-3.081050418e-07 pkt1=2.182606528e-13 kt2=4.671301857e-01 lkt2=-5.511902008e-07 wkt2=-3.249848058e-07 pkt2=3.588985769e-13 at=9.019482680e+03 lat=2.262838777e-01 wat=8.846774109e-02 pat=-1.917866080e-7 ute=1.741548466e+01 lute=-1.783883224e-05 wute=-1.199591092e-05 pute=1.158231248e-11 ua1=5.630177954e-08 lua1=-5.397351870e-14 wua1=-3.508084813e-14 pua1=3.440513481e-20 ub1=-4.245147974e-17 lub1=4.004881629e-23 wub1=2.631512563e-23 pub1=-2.524138019e-29 uc1=-1.081824386e-09 luc1=9.225882190e-16 wuc1=6.994086697e-16 puc1=-5.775545747e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.86 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='1.002349301e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.080230570e-07 wvth0=-2.800459028e-07 pvth0=1.333399360e-13 k1=-5.019757873e-01 lk1=4.651657491e-07 wk1=6.860620979e-07 pk1=-3.266588630e-13 k2=3.213237447e-01 lk2=-1.582948112e-07 wk2=-2.353313838e-07 pk2=1.120497438e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-3.779586465e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.115692428e-07 wvoff=1.526826335e-07 pvoff=-7.269769837e-14 nfactor=-1.116460866e+01 lnfactor=6.736309639e-06 wnfactor=8.456231739e-06 pnfactor=-4.026316355e-12 eta0=-4.616708363e-01 leta0=4.531247453e-07 weta0=-4.578546857e-13 peta0=2.180010989e-19 etab=-1.641277800e-01 letab=7.784955966e-8 u0=1.157814824e-02 lu0=5.434164814e-09 wu0=1.000406078e-08 pu0=-4.763293485e-15 ua=-4.719923498e-09 lua=1.556068250e-15 wua=2.358125433e-15 pua=-1.122788411e-21 ub=6.166566058e-18 lub=-2.033160645e-24 wub=-2.708631692e-24 pub=1.289677060e-30 uc=4.892255971e-10 luc=-2.079231619e-16 wuc=-2.801246538e-16 puc=1.333774322e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=8.467276777e+04 lvsat=4.849456217e-02 wvsat=-6.029030502e-02 pvsat=2.870638467e-8 a0=-7.247776846e+00 la0=4.110185382e-06 wa0=5.015157086e-06 pa0=-2.387896834e-12 ags=-6.434486981e+00 lags=3.138087144e-06 wags=5.290437637e-06 pags=-2.518967815e-12 a1=0.0 a2=0.42385546 b0=-1.501628594e-06 lb0=7.149794320e-13 wb0=1.045556960e-12 pb0=-4.978273089e-19 b1=-2.897519808e-08 lb1=1.379613491e-14 wb1=2.017490887e-14 pb1=-9.606000411e-21 keta=9.751614542e-01 lketa=-4.676963786e-07 wketa=-6.613034043e-07 pketa=3.148703577e-13 dwg=0.0 dwb=0.0 pclm=-1.480429790e+00 lpclm=9.200089246e-07 wpclm=1.666865769e-06 ppclm=-7.936547997e-13 pdiblc1=4.237879451e-01 lpdiblc1=-1.860530712e-07 wpdiblc1=1.434343351e-07 ppdiblc1=-6.829425058e-14 pdiblc2=2.591690982e-02 lpdiblc2=-1.231786313e-08 wpdiblc2=-1.018306457e-08 ppdiblc2=4.848523631e-15 pdiblcb=-6.530989907e-01 lpdiblcb=2.659189948e-07 wpdiblcb=4.503553757e-07 ppdiblcb=-2.144304072e-13 drout=-7.046982730e+00 ldrout=3.831458121e-06 wdrout=4.783699729e-06 pdrout=-2.277691654e-12 pscbe1=2.015071226e+09 lpscbe1=-7.514017517e+02 wpscbe1=-6.053099923e+02 ppscbe1=2.882098785e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-7.587468680e-05 lalpha0=3.798360027e-11 walpha0=5.028343301e-11 palpha0=-2.394175266e-17 alpha1=-1.460864150e+00 lalpha1=1.100285613e-06 walpha1=1.401035338e-06 palpha1=-6.670833619e-13 beta0=-3.749724754e+01 lbeta0=2.643280790e-05 wbeta0=3.300216575e-05 pbeta0=-1.571351919e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=1.554099991e-03 lkt1=-1.335579002e-07 wkt1=-1.649835406e-07 pkt1=7.855460309e-14 kt2=-1.554491249e-01 lkt2=5.653187723e-08 wkt2=8.333841687e-08 pkt2=-3.968042045e-14 at=4.600295332e+05 lat=-2.139632689e-01 wat=-2.108601223e-01 pat=1.003980952e-7 ute=-4.301595081e-01 lute=-4.190565268e-07 wute=-2.546560291e-07 pute=1.212509031e-13 ua1=1.177374702e-09 lua1=-1.646026586e-16 wua1=3.229120899e-16 pua1=-1.537500708e-22 ub1=-2.177482010e-18 lub1=7.359172347e-25 wub1=8.915225567e-25 pub1=-4.244859841e-31 uc1=-2.723054692e-10 luc1=1.323876614e-16 wuc1=2.103268131e-16 puc1=-1.001441675e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.87 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.094315479e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.094076978e-8 k1=8.414013965e-02 lk1=1.860948561e-7 k2=1.063879477e-01 lk2=-5.595614061e-08 wk2=1.387778781e-23 pk2=1.040834086e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425678e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663643e-8 nfactor=3.588363944e+00 lnfactor=-2.881117239e-07 wnfactor=3.552713679e-21 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=1.040834086e-23 petab=-1.301042607e-30 u0=1.975546521e-02 lu0=1.540649821e-9 ua=-1.703807103e-09 lua=1.199866544e-16 ub=1.993090002e-18 lub=-4.601845034e-26 uc=1.633443546e-11 luc=1.723734427e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.942043876e+05 lvsat=-3.657385172e-3 a0=1.280215623e+00 la0=4.970115974e-8 ags=-8.330949981e-01 lags=4.710627705e-07 pags=-5.551115123e-29 a1=0.0 a2=0.42385546 b0=3.484793983e-17 lb0=-7.880373722e-24 b1=-2.675520754e-18 lb1=6.050315613e-25 keta=6.166340678e-02 lketa=-3.274707228e-08 wketa=-1.387778781e-23 dwg=0.0 dwb=0.0 pclm=6.446949620e-01 lpclm=-9.183947440e-8 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 wpdiblc1=-5.551115123e-23 ppdiblc1=-2.775557562e-29 pdiblc2=-7.515255686e-03 lpdiblc2=3.600394425e-09 wpdiblc2=1.843143693e-24 ppdiblc2=3.117081246e-31 pdiblcb=-8.674421607e-02 lpdiblcb=-3.742902200e-9 drout=1.449262699e+00 ldrout=-2.139101923e-7 pscbe1=1.163107030e+08 lpscbe1=1.526664888e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183450e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126009e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532619e+03 lat=7.780439653e-3 ute=-1.302351205e+00 lute=-3.774660934e-9 ua1=1.605522255e-09 lua1=-3.684591219e-16 wua1=-8.271806126e-31 ub1=-1.843635241e-18 lub1=5.769607696e-25 wub1=7.703719778e-40 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=-1.292469707e-32 puc1=1.615587134e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.88 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820277676e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033728658e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217056813e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944838817e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083471173e-16 ags=1.250000000e+00 lags=4.460787295e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566857920e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563461134e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831734847e-18 drout=5.033266588e-01 ldrout=1.889157719e-16 pscbe1=7.914198799e+08 lpscbe1=1.866340637e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.132038907e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135939962e-25 ub1=7.077531681e-19 lub1=3.034206331e-34 uc1=1.471862500e-10 luc1=-4.393363028e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.89 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.5e-07 wmax=7.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='9.046558635e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.223929776e-08 wvth0=3.500080497e-07 pvth0=-5.464885685e-14 k1=0.90707349 k2=-2.212298632e-01 lk2=1.361869753e-08 wk2=4.273468679e-08 pk2=-6.672423057e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999998e-03 lcdscd=3.262303622e-19 wcdscd=2.012161271e-18 pcdscd=-3.141705646e-25 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749067557e-17 nfactor=4.984644527e+00 lnfactor=-3.918882146e-07 wnfactor=-1.521716776e-06 pnfactor=2.375947705e-13 eta0=1.166700699e-09 leta0=-1.471364695e-16 weta0=5.265131670e-19 peta0=-8.220765985e-26 etab=-0.043998 u0=8.366079997e-02 lu0=-8.526184836e-09 wu0=-3.121298300e-08 pu0=4.873470314e-15 ua=-1.167043358e-09 lua=-2.205575086e-18 wua=-8.564331521e-18 pua=1.337200466e-24 ub=-6.524880699e-20 lub=3.242009357e-25 wub=1.258884510e-24 pub=-1.965571919e-31 uc=7.700399986e-11 luc=1.717288990e-26 wuc=-1.381391623e-28 puc=2.155839471e-35 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.028209694e+05 lvsat=-2.614874881e-03 wvsat=6.045571396e-03 pvsat=-9.439313354e-10 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000007e-02 lketa=9.226508446e-18 wketa=7.893685705e-20 pketa=-1.232347557e-26 dwg=0.0 dwb=0.0 pclm=1.083066820e+00 lpclm=-1.411003228e-07 wpclm=-5.478978956e-07 ppclm=8.554658583e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.058713578e-24 walpha0=-1.577598864e-25 palpha0=2.463012992e-32 alpha1=0.85 beta0=1.057036139e+01 lbeta0=5.141203221e-07 wbeta0=1.996348684e-06 pbeta0=-3.117018981e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-6.697880826e-02 lkt1=-2.570601627e-08 wkt1=-9.981743435e-08 pkt1=1.558509493e-14 kt2=-0.028878939 at=5.372048692e+04 lat=1.012865687e-11 wat=-3.352761269e-14 pat=5.267793313e-21 ute=-2.138952857e+00 lute=1.285300811e-07 wute=4.990871718e-07 pute=-7.792547465e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.90 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.91 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-7 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-8 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 wub=-1.232595164e-38 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-7 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-7 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-07 wkt2=2.220446049e-22 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-6 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 puc1=3.308722450e-36 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.92 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-07 pk2=8.881784197e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 wua=-6.617444900e-30 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-8 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 wpclm=-8.881784197e-22 ppclm=1.065814104e-26 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-08 ppdiblc2=-5.551115123e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.93 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-8 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-6 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 pb1=-5.293955920e-35 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-8 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 ub1=-1.486104833e-18 lub1=3.235003467e-24 pub1=-1.232595164e-44 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.94 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-07 wnfactor=2.842170943e-20 eta0=-1.482776250e-03 leta0=3.918235528e-09 peta0=-6.938893904e-30 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=1.318389842e-22 petab=-3.538835891e-28 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 wuc=-4.135903063e-31 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-6 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 wketa=-5.551115123e-23 pketa=2.220446049e-28 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 walpha0=6.776263578e-27 palpha0=9.317362420e-33 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-7 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-02 wat=-9.313225746e-16 ute=-2.370540520e+00 lute=1.265004727e-6 ua1=-1.560482787e-09 lua1=2.774223792e-15 pua1=3.308722450e-36 ub1=9.526220239e-19 lub1=-1.584252469e-24 wub1=-3.081487911e-39 pub1=3.081487911e-45 uc1=7.177850760e-11 luc1=-3.002883819e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.95 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.404422957e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.190749679e-8 k1=6.296133048e-01 lk1=-7.362455486e-8 k2=-6.683124558e-02 lk2=2.651975321e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242963e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338157294e-9 nfactor=2.783078620e+00 lnfactor=9.531360915e-8 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=1.193489751e-21 peta0=5.412337245e-28 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.807882083e-02 lu0=-2.422399434e-9 ua=-8.304373629e-10 lua=-2.958561203e-16 ub=1.698955783e-18 lub=9.402944022e-26 uc=2.718870036e-11 luc=1.206923800e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.476990910e+04 lvsat=9.584280056e-2 a0=1.024210589e+00 la0=1.715943729e-7 ags=2.291547499e+00 lags=-1.016692010e-6 a1=0.0 a2=0.42385546 b0=2.229104169e-07 lb0=-1.061356743e-13 b1=4.301245672e-09 lb1=-2.047977910e-15 keta=-1.155907112e-01 lketa=5.164999443e-8 dwg=0.0 dwb=0.0 pclm=1.268894400e+00 lpclm=-3.890432982e-7 pdiblc1=6.603681753e-01 lpdiblc1=-2.986974357e-7 pdiblc2=9.120988834e-03 lpdiblc2=-4.320720496e-09 ppdiblc2=2.775557562e-29 pdiblcb=8.971602891e-02 lpdiblcb=-8.776197740e-08 wpdiblcb=1.647987302e-22 ppdiblcb=-2.203098814e-28 drout=8.432395257e-01 ldrout=7.463925758e-8 pscbe1=1.016674453e+09 lpscbe1=-2.760291058e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680640e-06 lalpha0=-1.505866109e-12 walpha0=5.421010862e-26 alpha1=0.85 beta0=1.693644131e+01 lbeta0=5.149690257e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693353e-01 lkt1=-3.990136186e-9 kt2=-1.799095058e-02 lkt2=-8.916908083e-9 at=1.122373799e+05 lat=-4.836690423e-2 ute=-8.501885195e-01 lute=-2.190655934e-7 ua1=1.709985088e-09 lua1=-4.181976372e-16 ub1=-7.070069559e-19 lub1=3.577112441e-26 uc1=7.460704527e-11 luc1=-3.278987563e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.96 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.094315479e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.094076978e-8 k1=8.414013965e-02 lk1=1.860948561e-7 k2=1.063879477e-01 lk2=-5.595614061e-08 wk2=2.220446049e-22 pk2=-8.326672685e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425678e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663643e-8 nfactor=3.588363944e+00 lnfactor=-2.881117239e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=-7.632783294e-23 petab=-4.510281038e-29 u0=1.975546521e-02 lu0=1.540649821e-9 ua=-1.703807103e-09 lua=1.199866544e-16 ub=1.993090002e-18 lub=-4.601845034e-26 uc=1.633443546e-11 luc=1.723734427e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.942043876e+05 lvsat=-3.657385172e-3 a0=1.280215623e+00 la0=4.970115974e-8 ags=-8.330949981e-01 lags=4.710627705e-07 wags=1.776356839e-21 pags=1.332267630e-27 a1=0.0 a2=0.42385546 b0=3.484793983e-17 lb0=-7.880373722e-24 b1=-2.675520754e-18 lb1=6.050315613e-25 keta=6.166340678e-02 lketa=-3.274707228e-08 wketa=1.665334537e-22 pketa=4.163336342e-29 dwg=0.0 dwb=0.0 pclm=6.446949620e-01 lpclm=-9.183947440e-08 wpclm=3.552713679e-21 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 wpdiblc1=-4.440892099e-22 ppdiblc1=-1.110223025e-28 pdiblc2=-7.515255686e-03 lpdiblc2=3.600394425e-09 wpdiblc2=4.336808690e-25 ppdiblc2=8.456776945e-30 pdiblcb=-8.674421607e-02 lpdiblcb=-3.742902200e-9 drout=1.449262699e+00 ldrout=-2.139101923e-7 pscbe1=1.163107030e+08 lpscbe1=1.526664888e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183450e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126009e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532619e+03 lat=7.780439653e-03 pat=-2.910383046e-23 ute=-1.302351205e+00 lute=-3.774660934e-9 ua1=1.605522255e-09 lua1=-3.684591219e-16 ub1=-1.843635241e-18 lub1=5.769607696e-25 wub1=6.162975822e-39 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=-2.584939414e-31 puc1=5.169878828e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.97 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820144449e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033839681e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217143549e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944977595e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083524464e-16 ags=1.250000000e+00 lags=4.461497838e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566924534e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.562906023e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831512802e-18 drout=5.033266588e-01 ldrout=1.889137735e-16 pscbe1=7.914198799e+08 lpscbe1=1.866149902e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.132094418e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135939574e-25 ub1=7.077531681e-19 lub1=3.034217886e-34 uc1=1.471862500e-10 luc1=-4.392329053e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.98 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.4e-07 wmax=6.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.030118625e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-7.090183690e-07 wvth0=-2.644814674e-06 pvth0=4.129507839e-13 k1=0.90707349 k2=-2.873543739e-01 lk2=2.394311414e-08 wk2=8.282478742e-08 pk2=-1.293193101e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.45863 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000024e-03 lcdscd=-3.677003146e-18 wcdscd=-1.353256396e-17 pcdscd=2.112914010e-24 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749178580e-17 nfactor=4.984644660e+00 lnfactor=-3.918882354e-07 wnfactor=-1.521716856e-06 pnfactor=2.375947830e-13 eta0=1.166700809e-09 leta0=-1.471364686e-16 weta0=5.265167660e-19 peta0=-8.220822178e-26 etab=-0.043998 u0=-2.244160702e-01 lu0=3.957570537e-08 wu0=1.555684780e-07 pu0=-2.428983988e-14 ua=-1.167043295e-09 lua=-2.205584809e-18 wua=-8.564369276e-18 pua=1.337206361e-24 ub=-6.524872088e-20 lub=3.242009223e-25 wub=1.258884458e-24 pub=-1.965571837e-31 uc=7.700399986e-11 luc=1.744689348e-26 wuc=9.280966473e-28 puc=-1.449634023e-34 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.450773213e+06 lvsat=2.555707064e-01 wvsat=1.008589960e+00 pvsat=-1.574772019e-7 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000007e-02 lketa=9.068967799e-18 wketa=-5.320188734e-19 pketa=8.304468224e-26 dwg=0.0 dwb=0.0 pclm=1.083066832e+00 lpclm=-1.411003247e-07 wpclm=-5.478979030e-07 ppclm=8.554658699e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000001e-08 lalpha0=-1.744040838e-24 walpha0=1.064720415e-24 palpha0=-1.662302159e-31 alpha1=0.85 beta0=1.057036138e+01 lbeta0=5.141203238e-07 wbeta0=1.996348691e-06 pbeta0=-3.117018992e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-6.697881003e-02 lkt1=-2.570601599e-08 wkt1=-9.981743328e-08 pkt1=1.558509476e-14 kt2=-0.028878939 at=5.372048692e+04 lat=1.019611955e-11 wat=2.272427082e-13 pat=-3.562308848e-20 ute=-2.138952848e+00 lute=1.285300797e-07 wute=4.990871664e-07 pute=-7.792547381e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.99 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.100 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-7 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-8 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-7 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 wb0=-5.293955920e-29 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-07 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-7 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-6 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.101 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-07 pk2=-2.220446049e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-8 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 wpclm=2.220446049e-22 ppclm=-5.329070518e-27 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-08 ppdiblc2=-2.775557562e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 wua1=-3.308722450e-30 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 wuc1=5.169878828e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.102 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-8 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-06 wa0=3.552713679e-21 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-8 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 ub1=-1.486104833e-18 lub1=3.235003467e-24 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.103 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-7 eta0=-1.482776250e-03 leta0=3.918235528e-09 peta0=-1.734723476e-30 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=-3.122502257e-23 petab=-3.989863995e-29 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-06 pags=1.776356839e-27 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 wketa=-2.775557562e-23 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 walpha0=2.646977960e-27 palpha0=5.505714157e-33 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-07 wkt1=8.881784197e-22 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-2 ute=-2.370540520e+00 lute=1.265004727e-6 ua1=-1.560482787e-09 lua1=2.774223792e-15 wua1=1.240770919e-30 pua1=3.308722450e-36 ub1=9.526220239e-19 lub1=-1.584252469e-24 wub1=-3.851859889e-40 pub1=7.703719778e-46 uc1=7.177850760e-11 luc1=-3.002883819e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.104 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.404422957e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.190749679e-8 k1=6.296133048e-01 lk1=-7.362455486e-8 k2=-6.683124558e-02 lk2=2.651975321e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242963e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338157294e-9 nfactor=2.783078620e+00 lnfactor=9.531360915e-8 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=4.232725281e-22 peta0=2.081668171e-29 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.807882083e-02 lu0=-2.422399434e-9 ua=-8.304373629e-10 lua=-2.958561203e-16 ub=1.698955783e-18 lub=9.402944022e-26 uc=2.718870036e-11 luc=1.206923800e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.476990910e+04 lvsat=9.584280056e-2 a0=1.024210589e+00 la0=1.715943729e-7 ags=2.291547499e+00 lags=-1.016692010e-6 a1=0.0 a2=0.42385546 b0=2.229104169e-07 lb0=-1.061356743e-13 b1=4.301245672e-09 lb1=-2.047977910e-15 keta=-1.155907112e-01 lketa=5.164999443e-8 dwg=0.0 dwb=0.0 pclm=1.268894400e+00 lpclm=-3.890432982e-7 pdiblc1=6.603681753e-01 lpdiblc1=-2.986974357e-7 pdiblc2=9.120988834e-03 lpdiblc2=-4.320720496e-9 pdiblcb=8.971602891e-02 lpdiblcb=-8.776197740e-08 wpdiblcb=4.770489559e-23 ppdiblcb=-1.951563910e-29 drout=8.432395257e-01 ldrout=7.463925758e-8 pscbe1=1.016674453e+09 lpscbe1=-2.760291058e+02 wpscbe1=-1.907348633e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680640e-06 lalpha0=-1.505866109e-12 walpha0=-1.355252716e-26 alpha1=0.85 beta0=1.693644131e+01 lbeta0=5.149690257e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693353e-01 lkt1=-3.990136186e-9 kt2=-1.799095058e-02 lkt2=-8.916908083e-9 at=1.122373799e+05 lat=-4.836690423e-2 ute=-8.501885195e-01 lute=-2.190655934e-7 ua1=1.709985088e-09 lua1=-4.181976372e-16 ub1=-7.070069559e-19 lub1=3.577112441e-26 uc1=7.460704527e-11 luc1=-3.278987563e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.105 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.094315479e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.094076978e-8 k1=8.414013965e-02 lk1=1.860948561e-7 k2=1.063879477e-01 lk2=-5.595614061e-08 wk2=5.551115123e-23 pk2=4.857225733e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425678e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663643e-8 nfactor=3.588363944e+00 lnfactor=-2.881117239e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=-3.469446952e-24 petab=-3.035766083e-30 u0=1.975546521e-02 lu0=1.540649821e-9 ua=-1.703807103e-09 lua=1.199866544e-16 ub=1.993090002e-18 lub=-4.601845034e-26 uc=1.633443546e-11 luc=1.723734427e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.942043876e+05 lvsat=-3.657385172e-03 wvsat=-4.656612873e-16 a0=1.280215623e+00 la0=4.970115974e-8 ags=-8.330949981e-01 lags=4.710627705e-07 wags=-8.881784197e-22 pags=1.110223025e-28 a1=0.0 a2=0.42385546 b0=3.484793983e-17 lb0=-7.880373722e-24 b1=-2.675520754e-18 lb1=6.050315613e-25 keta=6.166340678e-02 lketa=-3.274707228e-08 wketa=2.775557562e-23 pketa=-2.081668171e-29 dwg=0.0 dwb=0.0 pclm=6.446949620e-01 lpclm=-9.183947440e-8 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 ppdiblc1=-1.110223025e-28 pdiblc2=-7.515255686e-03 lpdiblc2=3.600394425e-09 wpdiblc2=1.734723476e-24 ppdiblc2=-4.878909776e-31 pdiblcb=-8.674421607e-02 lpdiblcb=-3.742902200e-9 drout=1.449262699e+00 ldrout=-2.139101923e-7 pscbe1=1.163107030e+08 lpscbe1=1.526664888e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183450e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126009e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532619e+03 lat=7.780439653e-03 pat=7.275957614e-24 ute=-1.302351205e+00 lute=-3.774660934e-9 ua1=1.605522255e-09 lua1=-3.684591219e-16 ub1=-1.843635241e-18 lub1=5.769607696e-25 pub1=3.851859889e-46 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=-1.033975766e-31 puc1=4.523643975e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.106 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820144449e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033750863e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217074161e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944811062e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083488937e-16 ags=1.250000000e+00 lags=4.460964931e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566880125e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563599912e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831734847e-18 drout=5.033266588e-01 ldrout=1.889164380e-16 pscbe1=7.914198799e+08 lpscbe1=1.866340637e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.132038907e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135939574e-25 ub1=7.077531681e-19 lub1=3.034202479e-34 uc1=1.471862500e-10 luc1=-4.393156233e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.107 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.1e-07 wmax=6.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='-1.524716387e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.144273503e-07 wvth0=1.263715457e-06 pvth0=-1.973114765e-13 k1=0.90707349 k2=-1.638207879e-01 lk2=4.655074161e-09 wk2=9.163933717e-09 pk2=-1.430819955e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585131626e-01 ldsub=1.824252398e-11 wdsub=6.966803737e-11 pdsub=-1.087768868e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.335147271e-19 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749045353e-17 nfactor=6.350352411e+00 lnfactor=-6.051243808e-07 wnfactor=-2.336063805e-06 pnfactor=3.647436583e-13 eta0=1.641780072e-02 leta0=-2.563409442e-09 weta0=-9.789637375e-09 peta0=1.528514821e-15 etab=-0.043998 u0=-4.312098015e-02 lu0=1.126901519e-08 wu0=4.746547912e-08 pu0=-7.411070048e-15 ua=-1.067214444e-09 lua=-1.779246228e-17 wua=-6.809051619e-17 pua=1.063138084e-23 ub=7.948211664e-18 lub=-9.269887284e-25 wub=-3.519397727e-24 pub=5.495046835e-31 uc=3.253499464e-10 luc=-3.877574270e-17 wuc=-1.480842177e-16 puc=2.312127742e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.172496790e+06 lvsat=-1.540161788e-01 wvsat=-5.556187243e-01 pvsat=8.675208514e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000007e-02 lketa=9.208467322e-18 dwg=0.0 dwb=0.0 pclm=-2.993692896e-01 lpclm=7.474772162e-08 wpclm=2.764238727e-07 ppclm=-4.315971778e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.022661738e-24 alpha1=0.85 beta0=1.391835560e+01 lbeta0=-8.622102004e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.708984644e-01 lkt1=3.736038317e-08 wkt1=1.410325861e-07 pkt1=-2.202026386e-14 kt2=-0.028878939 at=5.372048692e+04 lat=1.013639849e-11 ute=2.117733343e-01 lute=-2.385029035e-07 wute=-9.026085430e-07 pute=1.409296875e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.108 nmos lmin=2.0e-05 lmax=0.0001 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.109 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-7 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-8 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-7 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-7 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-07 wkt2=2.220446049e-22 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-06 wute=7.105427358e-21 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.110 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-07 pk2=-4.440892099e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 wua=-6.617444900e-30 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-08 wketa=-5.551115123e-23 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 wpclm=-8.881784197e-22 ppclm=5.329070518e-27 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 wuc1=-2.067951531e-31 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.111 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-8 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-6 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 pb1=5.293955920e-35 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-8 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 ub1=-1.486104833e-18 lub1=3.235003467e-24 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.112 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-7 eta0=-1.482776250e-03 leta0=3.918235528e-09 peta0=-6.938893904e-30 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=1.387778781e-23 petab=-2.081668171e-29 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 pua=-3.308722450e-36 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-6 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 walpha0=7.623296525e-27 palpha0=-2.159934015e-32 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-7 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-2 ute=-2.370540520e+00 lute=1.265004727e-06 wute=1.421085472e-20 ua1=-1.560482787e-09 lua1=2.774223792e-15 wua1=1.654361225e-30 pua1=-4.963083675e-36 ub1=9.526220239e-19 lub1=-1.584252469e-24 wub1=1.540743956e-39 pub1=1.540743956e-45 uc1=7.177850760e-11 luc1=-3.002883819e-17 wuc1=4.135903063e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.113 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.404422957e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.190749679e-8 k1=6.296133048e-01 lk1=-7.362455486e-8 k2=-6.683124558e-02 lk2=2.651975321e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242963e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338157294e-9 nfactor=2.783078620e+00 lnfactor=9.531360915e-8 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=3.885780586e-22 peta0=-3.885780586e-28 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.807882083e-02 lu0=-2.422399434e-9 ua=-8.304373629e-10 lua=-2.958561203e-16 ub=1.698955783e-18 lub=9.402944022e-26 uc=2.718870036e-11 luc=1.206923800e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-1.476990910e+04 lvsat=9.584280056e-2 a0=1.024210589e+00 la0=1.715943729e-7 ags=2.291547499e+00 lags=-1.016692010e-6 a1=0.0 a2=0.42385546 b0=2.229104169e-07 lb0=-1.061356743e-13 b1=4.301245672e-09 lb1=-2.047977910e-15 keta=-1.155907112e-01 lketa=5.164999443e-8 dwg=0.0 dwb=0.0 pclm=1.268894400e+00 lpclm=-3.890432982e-7 pdiblc1=6.603681753e-01 lpdiblc1=-2.986974357e-7 pdiblc2=9.120988834e-03 lpdiblc2=-4.320720496e-9 pdiblcb=8.971602891e-02 lpdiblcb=-8.776197740e-08 wpdiblcb=6.765421556e-23 ppdiblcb=7.632783294e-29 drout=8.432395257e-01 ldrout=7.463925758e-8 pscbe1=1.016674453e+09 lpscbe1=-2.760291058e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680640e-06 lalpha0=-1.505866109e-12 alpha1=0.85 beta0=1.693644131e+01 lbeta0=5.149690257e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693353e-01 lkt1=-3.990136186e-9 kt2=-1.799095058e-02 lkt2=-8.916908083e-9 at=1.122373799e+05 lat=-4.836690423e-2 ute=-8.501885195e-01 lute=-2.190655934e-7 ua1=1.709985088e-09 lua1=-4.181976372e-16 ub1=-7.070069559e-19 lub1=3.577112441e-26 uc1=7.460704527e-11 luc1=-3.278987563e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.114 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.094315479e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.094076978e-8 k1=8.414013965e-02 lk1=1.860948561e-7 k2=1.063879477e-01 lk2=-5.595614061e-08 wk2=-2.220446049e-22 pk2=-5.551115123e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425678e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663643e-8 nfactor=3.588363944e+00 lnfactor=-2.881117239e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=6.245004514e-23 petab=5.204170428e-30 u0=1.975546521e-02 lu0=1.540649821e-9 ua=-1.703807103e-09 lua=1.199866544e-16 ub=1.993090002e-18 lub=-4.601845034e-26 uc=1.633443546e-11 luc=1.723734427e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.942043876e+05 lvsat=-3.657385172e-3 a0=1.280215623e+00 la0=4.970115974e-8 ags=-8.330949981e-01 lags=4.710627705e-07 pags=4.440892099e-28 a1=0.0 a2=0.42385546 b0=3.484793983e-17 lb0=-7.880373722e-24 b1=-2.675520754e-18 lb1=6.050315613e-25 keta=6.166340678e-02 lketa=-3.274707228e-08 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=6.446949620e-01 lpclm=-9.183947440e-8 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 ppdiblc1=1.110223025e-28 pdiblc2=-7.515255686e-03 lpdiblc2=3.600394425e-09 wpdiblc2=1.214306433e-23 ppdiblc2=-3.252606517e-31 pdiblcb=-8.674421607e-02 lpdiblcb=-3.742902200e-9 drout=1.449262699e+00 ldrout=-2.139101923e-7 pscbe1=1.163107030e+08 lpscbe1=1.526664888e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183450e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126009e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532619e+03 lat=7.780439653e-3 ute=-1.302351205e+00 lute=-3.774660934e-9 ua1=1.605522255e-09 lua1=-3.684591219e-16 ub1=-1.843635241e-18 lub1=5.769607696e-25 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=1.550963649e-31 puc1=-2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.115 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820499721e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033662045e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217074161e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944977595e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083453410e-16 ags=1.250000000e+00 lags=4.460787295e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.567102169e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563461134e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831512802e-18 drout=5.033266588e-01 ldrout=1.889155499e-16 pscbe1=7.914198799e+08 lpscbe1=1.866531372e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.131983396e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135940608e-25 ub1=7.077531681e-19 lub1=3.034217886e-34 uc1=1.471862500e-10 luc1=-4.393156233e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.116 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=6.0e-07 wmax=6.1e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='2.866190766e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.161267641e-08 wvth0=2.379887877e-07 pvth0=-3.715861736e-14 k1=0.90707349 k2=-1.315305804e-01 lk2=-3.865896863e-10 wk2=-9.121429602e-09 pk2=1.424183532e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585131590e-01 ldsub=1.824309235e-11 wdsub=6.967009877e-11 pdsub=-1.087801054e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.335043187e-19 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749089762e-17 nfactor=6.350352394e+00 lnfactor=-6.051243782e-07 wnfactor=-2.336063796e-06 pnfactor=3.647436568e-13 eta0=1.641776644e-02 leta0=-2.563404346e-09 weta0=-9.789618892e-09 peta0=1.528511935e-15 etab=-0.043998 u0=-1.256786806e-01 lu0=2.415924431e-08 wu0=9.421641885e-08 pu0=-1.471057477e-14 ua=-1.067214413e-09 lua=-1.779246712e-17 wua=-6.809053374e-17 pua=1.063138358e-23 ub=7.948211668e-18 lub=-9.269887290e-25 wub=-3.519397730e-24 pub=5.495046839e-31 uc=3.253499468e-10 luc=-3.877574275e-17 wuc=-1.480842179e-16 puc=2.312127745e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.813028449e+05 lvsat=7.448790184e-04 wvsat=5.676565231e-03 pvsat=-8.863161888e-10 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000007e-02 lketa=9.208189766e-18 dwg=0.0 dwb=0.0 pclm=-2.993692910e-01 lpclm=7.474772183e-08 wpclm=2.764238734e-07 ppclm=-4.315971790e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.022714678e-24 alpha1=0.85 beta0=1.391835560e+01 lbeta0=-8.622102004e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.708984687e-01 lkt1=3.736038383e-08 wkt1=1.410325885e-07 pkt1=-2.202026424e-14 kt2=-0.028878939 at=5.372048692e+04 lat=1.013628207e-11 ute=2.117733753e-01 lute=-2.385029099e-07 wute=-9.026085663e-07 pute=1.409296911e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.117 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.118 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-07 wk1=-1.776356839e-21 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-8 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-7 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-07 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+03 ppscbe1=-7.629394531e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-7 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-6 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 wuc1=1.033975766e-31 puc1=8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.119 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-07 pk2=2.220446049e-28 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-08 wketa=-2.775557562e-23 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 wuc1=-1.033975766e-31 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.120 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-08 wvoff=-4.440892099e-22 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-6 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-08 wpdiblcb=-1.110223025e-22 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 ub1=-1.486104833e-18 lub1=3.235003467e-24 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.121 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-7 eta0=-1.482776250e-03 leta0=3.918235528e-09 weta0=1.734723476e-24 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=-7.112366252e-23 petab=-1.457167720e-28 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-6 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 pketa=-8.326672685e-29 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 walpha0=-5.082197684e-27 palpha0=-4.658681210e-33 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-7 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-2 ute=-2.370540520e+00 lute=1.265004727e-06 wute=7.105427358e-21 ua1=-1.560482787e-09 lua1=2.774223792e-15 wua1=8.271806126e-31 pua1=-1.654361225e-36 ub1=9.526220239e-19 lub1=-1.584252469e-24 pub1=7.703719778e-46 uc1=7.177850760e-11 luc1=-3.002883819e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.122 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.069106764e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-5.297468249e-08 wvth0=-3.697516376e-08 pvth0=3.609278846e-14 k1=6.296133055e-01 lk1=-7.362455560e-08 wk1=-4.224496308e-16 pk1=4.123679176e-22 k2=-2.607336961e-02 lk2=-1.326547680e-08 wk2=-2.267287276e-08 pk2=2.213180732e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939289e-01 ldsub=4.676284059e-08 wdsub=-1.245989978e-16 pdsub=1.216262646e-22 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242954e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338158196e-09 wvoff=-5.140243786e-16 pvoff=5.017577465e-22 nfactor=2.783078629e+00 lnfactor=9.531360038e-08 wnfactor=-4.994376468e-15 pnfactor=4.875175819e-21 eta0=-4.616715920e-01 leta0=4.531251054e-07 weta0=2.850791964e-16 peta0=-2.782767558e-22 etab=-1.641277801e-01 letab=7.784955976e-08 wetab=5.727862629e-17 petab=-5.591149765e-23 u0=-1.160916747e-02 lu0=3.631847472e-08 wu0=2.207771351e-08 pu0=-2.155085096e-14 ua=-8.304373597e-10 lua=-2.958561234e-16 wua=-1.795418681e-24 pua=1.752574034e-30 ub=1.698955786e-18 lub=9.402943746e-26 wub=-1.572551074e-33 pub=1.535024714e-39 uc=2.718870047e-11 luc=1.206923788e-17 wuc=-6.421196300e-26 puc=6.267950752e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-3.875453975e+05 lvsat=4.597223747e-01 wvsat=2.073682942e-01 pvsat=-2.024196572e-7 a0=1.024210583e+00 la0=1.715943783e-07 wa0=3.105625979e-15 pa0=-3.031509266e-21 ags=2.291547474e+00 lags=-1.016691985e-06 wags=1.372291081e-14 pags=-1.339542877e-20 a1=0.0 a2=0.42385546 b0=2.229104165e-07 lb0=-1.061356738e-13 wb0=2.598993544e-22 pb0=-2.536971674e-28 b1=4.301245708e-09 lb1=-2.047977945e-15 wb1=-1.995430953e-23 pb1=1.947811157e-29 keta=-1.155907120e-01 lketa=5.164999526e-08 wketa=4.734999060e-16 pketa=-4.622001670e-22 dwg=0.0 dwb=0.0 pclm=1.268894407e+00 lpclm=-3.890433046e-07 wpclm=-3.627615541e-15 ppclm=3.541048343e-21 pdiblc1=6.603681741e-01 lpdiblc1=-2.986974345e-07 wpdiblc1=6.799645291e-16 ppdiblc1=-6.637375094e-22 pdiblc2=9.120988864e-03 lpdiblc2=-4.320720524e-09 wpdiblc2=-1.638658653e-17 ppdiblc2=1.599552435e-23 pdiblcb=8.971602867e-02 lpdiblcb=-8.776197717e-08 wpdiblcb=1.316537825e-16 ppdiblcb=-1.285117945e-22 drout=8.432395265e-01 ldrout=7.463925678e-08 wdrout=-4.569820078e-16 pdrout=4.460751768e-22 pscbe1=1.016674444e+09 lpscbe1=-2.760290966e+02 wpscbe1=5.261962891e-06 ppscbe1=-5.136388779e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680628e-06 lalpha0=-1.505866098e-12 walpha0=6.176455831e-21 palpha0=-6.029058546e-27 alpha1=0.85 beta0=1.693644136e+01 lbeta0=5.149689774e-07 wbeta0=-2.750090289e-14 pbeta0=2.684464562e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693354e-01 lkt1=-3.990136108e-09 wkt1=4.413180932e-17 pkt1=-4.307931789e-23 kt2=-1.799095059e-02 lkt2=-8.916908071e-09 wkt2=7.193023954e-18 pkt2=-7.021383475e-24 at=1.122373789e+05 lat=-4.836690327e-02 wat=5.465282593e-10 pat=-5.334857851e-16 ute=-8.501885175e-01 lute=-2.190655954e-07 wute=-1.129670579e-15 pute=1.102709035e-21 ua1=1.709985083e-09 lua1=-4.181976331e-16 wua1=2.340299094e-24 pua1=-2.284447859e-30 ub1=-7.070069568e-19 lub1=3.577112531e-26 wub1=5.134590861e-34 pub1=-5.012040087e-40 uc1=7.460704537e-11 luc1=-3.278987573e-17 wuc1=-5.686804673e-26 puc1=5.551085014e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.123 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.764947864e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=9.121017709e-09 wvth0=7.395032753e-08 pvth0=-1.672283127e-14 k1=8.414013813e-02 lk1=1.860948564e-07 wk1=8.448974853e-16 pk1=-1.910622771e-22 k2=2.487219580e-02 lk2=-3.752249453e-08 wk2=4.534574552e-08 pk2=-1.025430551e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425674e-01 ldsub=6.388057806e-08 wdsub=2.491997719e-16 pdsub=-5.635314437e-23 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188898e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663601e-08 wvoff=1.028048757e-15 pvoff=-2.324788140e-22 nfactor=3.588363926e+00 lnfactor=-2.881117199e-07 wnfactor=9.988738725e-15 pnfactor=-2.258811804e-21 eta0=9.325986808e-01 leta0=-2.107371652e-07 weta0=-5.701608075e-16 peta0=1.289333085e-22 etab=3.860778713e-02 letab=-1.868014228e-08 wetab=-1.145570479e-16 petab=2.590545660e-23 u0=9.913144182e-02 lu0=-1.640911603e-08 wu0=-4.415542702e-08 pu0=9.985131645e-15 ua=-1.703807110e-09 lua=1.199866558e-16 wua=3.590843979e-24 pua=-8.120200463e-31 ub=1.993089997e-18 lub=-4.601844906e-26 wub=3.145102147e-33 pub=-7.112212766e-40 uc=1.633443523e-11 luc=1.723734432e-17 wuc=1.284239260e-25 puc=-2.904122563e-32 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.397553643e+05 lvsat=-1.722533008e-01 wvsat=-4.147365884e-01 pvsat=9.378687316e-8 a0=1.280215634e+00 la0=4.970115722e-08 wa0=-6.211244852e-15 pa0=1.404586669e-21 ags=-8.330949487e-01 lags=4.710627593e-07 wags=-2.744582339e-14 pags=6.206488878e-21 a1=0.0 a2=0.42385546 b0=9.692640833e-16 lb0=-2.191855027e-22 wb0=-5.197988811e-22 pb0=1.175452398e-28 b1=-7.441720181e-17 lb1=1.682840835e-23 wb1=3.990860582e-23 pb1=-9.024772486e-30 keta=6.166340848e-02 lketa=-3.274707267e-08 wketa=-9.469993401e-16 pketa=2.141506625e-22 dwg=0.0 dwb=0.0 pclm=6.446949490e-01 lpclm=-9.183947145e-08 wpclm=7.255232859e-15 ppclm=-1.640669378e-21 pdiblc1=-2.599865108e-01 lpdiblc1=1.395165637e-07 wpdiblc1=-1.359929169e-15 ppdiblc1=3.075291410e-22 pdiblc2=-7.515255745e-03 lpdiblc2=3.600394438e-09 wpdiblc2=3.277315311e-17 ppdiblc2=-7.411186628e-24 pdiblcb=-8.674421560e-02 lpdiblcb=-3.742902307e-09 wpdiblcb=-2.633075979e-16 ppdiblcb=5.954337023e-23 drout=1.449262698e+00 ldrout=-2.139101919e-07 wdrout=9.139604629e-16 pdrout=-2.066791183e-22 pscbe1=1.163107219e+08 lpscbe1=1.526664846e+02 wpscbe1=-1.052392387e-05 ppscbe1=2.379837990e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183472e-06 lalpha0=-1.670372440e-12 walpha0=-1.235289811e-20 palpha0=2.793436733e-27 alpha1=0.85 beta0=2.136300361e+01 lbeta0=-1.592676664e-06 wbeta0=5.500186262e-14 pbeta0=-1.243789427e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121571e-01 lkt1=1.636126006e-08 wkt1=-8.826450681e-17 pkt1=1.995958954e-23 kt2=-4.380991829e-02 lkt2=3.376431932e-09 wkt2=-1.438626995e-17 pkt2=3.253203262e-24 at=-5.685530654e+03 lat=7.780439208e-03 wat=-1.093056344e-09 pat=2.471793850e-16 ute=-1.302351209e+00 lute=-3.774660016e-09 wute=2.259334053e-15 pute=-5.109175305e-22 ua1=1.605522263e-09 lua1=-3.684591238e-16 wua1=-4.680594879e-24 pua1=1.058450386e-30 ub1=-1.843635239e-18 lub1=5.769607691e-25 wub1=-1.026915091e-33 pub1=2.322232401e-40 uc1=-1.222035416e-10 luc1=6.091872993e-17 wuc1=1.137358867e-25 puc1=-2.571980467e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.124 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820322085e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033750863e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217039466e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944755551e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083453410e-16 ags=1.250000000e+00 lags=4.460787295e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566835716e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563461134e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831734847e-18 drout=5.033266588e-01 ldrout=1.889155499e-16 pscbe1=7.914198799e+08 lpscbe1=1.866531372e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.132038907e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135940608e-25 ub1=7.077531681e-19 lub1=3.034217886e-34 uc1=1.471862500e-10 luc1=-4.393569824e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.125 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.8e-07 wmax=6.0e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='3.235046079e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.585351709e-08 wvth0=2.174700306e-07 pvth0=-3.395490070e-14 k1=0.90707349 k2=-4.369331416e-01 lk2=4.729774462e-08 wk2=1.607685180e-07 pk2=-2.510175332e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585131590e-01 ldsub=1.824309234e-11 wdsub=6.967009872e-11 pdsub=-1.087801053e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.335112576e-19 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749089762e-17 nfactor=6.350352394e+00 lnfactor=-6.051243782e-07 wnfactor=-2.336063796e-06 pnfactor=3.647436568e-13 eta0=1.641776644e-02 leta0=-2.563404346e-09 weta0=-9.789618892e-09 peta0=1.528511935e-15 etab=-0.043998 u0=2.566536566e-01 lu0=-3.553659750e-08 wu0=-1.184681784e-07 pu0=1.849714750e-14 ua=-1.067214413e-09 lua=-1.779246712e-17 wua=-6.809053374e-17 pua=1.063138358e-23 ub=7.948211668e-18 lub=-9.269887290e-25 wub=-3.519397730e-24 pub=5.495046839e-31 uc=3.253499468e-10 luc=-3.877574275e-17 wuc=-1.480842179e-16 puc=2.312127745e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.328009575e+05 lvsat=-7.295830301e-03 wvsat=-2.297090788e-02 pvsat=3.586585673e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000007e-02 lketa=9.208467322e-18 dwg=0.0 dwb=0.0 pclm=-2.993692910e-01 lpclm=7.474772183e-08 wpclm=2.764238734e-07 ppclm=-4.315971790e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.022608799e-24 alpha1=0.85 beta0=1.391835560e+01 lbeta0=-8.622102004e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.708984687e-01 lkt1=3.736038383e-08 wkt1=1.410325885e-07 pkt1=-2.202026424e-14 kt2=-0.028878939 at=5.372048692e+04 lat=1.013628207e-11 ute=2.117733753e-01 lute=-2.385029099e-07 wute=-9.026085663e-07 pute=1.409296911e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.126 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.127 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-7 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-8 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-7 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-07 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-7 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-6 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.128 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-8 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 wpclm=4.440892099e-22 ppclm=-8.881784197e-28 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 puc1=-4.135903063e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.129 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-8 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-6 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-8 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 ub1=-1.486104833e-18 lub1=3.235003467e-24 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.130 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-7 eta0=-1.482776250e-03 leta0=3.918235528e-9 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=4.683753385e-23 petab=8.326672685e-29 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 pua=-8.271806126e-37 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-6 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 pketa=8.326672685e-29 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 walpha0=7.411538288e-28 palpha0=6.140988868e-33 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-7 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-02 wat=2.328306437e-16 ute=-2.370540520e+00 lute=1.265004727e-6 ua1=-1.560482787e-09 lua1=2.774223792e-15 wua1=4.135903063e-31 pua1=8.271806126e-37 ub1=9.526220239e-19 lub1=-1.584252469e-24 wub1=-7.703719778e-40 pub1=-1.155557967e-45 uc1=7.177850760e-11 luc1=-3.002883819e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.131 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.379634364e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.432720057e-8 k1=6.296133047e-01 lk1=-7.362455483e-8 k2=-6.835126213e-02 lk2=2.800349610e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242964e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338157261e-9 nfactor=2.783078619e+00 lnfactor=9.531360947e-8 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=-4.163336342e-23 peta0=-3.295974604e-28 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.955893720e-02 lu0=-3.867194305e-9 ua=-8.304373631e-10 lua=-2.958561202e-16 ub=1.698955783e-18 lub=9.402944032e-26 uc=2.718870035e-11 luc=1.206923800e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-8.676901760e+02 lvsat=8.227234419e-2 a0=1.024210589e+00 la0=1.715943727e-7 ags=2.291547500e+00 lags=-1.016692010e-6 a1=0.0 a2=0.42385546 b0=2.229104170e-07 lb0=-1.061356743e-13 b1=4.301245670e-09 lb1=-2.047977909e-15 keta=-1.155907111e-01 lketa=5.164999439e-8 dwg=0.0 dwb=0.0 pclm=1.268894400e+00 lpclm=-3.890432980e-7 pdiblc1=6.603681753e-01 lpdiblc1=-2.986974357e-7 pdiblc2=9.120988833e-03 lpdiblc2=-4.320720495e-9 pdiblcb=8.971602892e-02 lpdiblcb=-8.776197741e-08 wpdiblcb=-5.377642776e-23 ppdiblcb=4.553649124e-30 drout=8.432395256e-01 ldrout=7.463925761e-8 pscbe1=1.016674454e+09 lpscbe1=-2.760291061e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680640e-06 lalpha0=-1.505866109e-12 alpha1=0.85 beta0=1.693644131e+01 lbeta0=5.149690275e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693353e-01 lkt1=-3.990136189e-9 kt2=-1.799095058e-02 lkt2=-8.916908084e-9 at=1.122373800e+05 lat=-4.836690427e-2 ute=-8.501885196e-01 lute=-2.190655934e-7 ua1=1.709985088e-09 lua1=-4.181976374e-16 ub1=-7.070069558e-19 lub1=3.577112438e-26 uc1=7.460704526e-11 luc1=-3.278987563e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.132 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.143892664e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.206188842e-8 k1=8.414013971e-02 lk1=1.860948561e-7 k2=1.094279808e-01 lk2=-5.664360154e-08 wk2=2.775557562e-23 pk2=-6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425679e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663645e-8 nfactor=3.588363944e+00 lnfactor=-2.881117241e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=-6.938893904e-24 petab=-7.372574773e-30 u0=1.679523247e-02 lu0=2.210065012e-9 ua=-1.703807103e-09 lua=1.199866543e-16 ub=1.993090003e-18 lub=-4.601845039e-26 uc=1.633443547e-11 luc=1.723734426e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.663999498e+05 lvsat=2.630199184e-3 a0=1.280215623e+00 la0=4.970115984e-8 ags=-8.330949999e-01 lags=4.710627709e-07 wags=4.440892099e-22 pags=4.440892099e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.166340672e-02 lketa=-3.274707227e-08 wketa=1.387778781e-23 pketa=2.775557562e-29 dwg=0.0 dwb=0.0 pclm=6.446949625e-01 lpclm=-9.183947451e-8 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 ppdiblc1=-1.110223025e-28 pdiblc2=-7.515255684e-03 lpdiblc2=3.600394425e-09 wpdiblc2=4.119968255e-24 ppdiblc2=-2.927345866e-30 pdiblcb=-8.674421609e-02 lpdiblcb=-3.742902196e-9 drout=1.449262700e+00 ldrout=-2.139101923e-7 pscbe1=1.163107023e+08 lpscbe1=1.526664890e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183449e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126010e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532692e+03 lat=7.780439669e-03 pat=7.275957614e-24 ute=-1.302351205e+00 lute=-3.774660968e-9 ua1=1.605522255e-09 lua1=-3.684591218e-16 ub1=-1.843635241e-18 lub1=5.769607696e-25 wub1=1.540743956e-39 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=1.292469707e-32 puc1=4.846761402e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.133 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820144449e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033750863e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217039466e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944811062e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083453410e-16 ags=1.250000000e+00 lags=4.460964931e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566880125e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563599912e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831734847e-18 drout=5.033266588e-01 ldrout=1.889155499e-16 pscbe1=7.914198799e+08 lpscbe1=1.866245270e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.132038907e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135939832e-25 ub1=7.077531681e-19 lub1=3.034202479e-34 uc1=1.471862500e-10 luc1=-4.393569824e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.134 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.5e-07 wmax=5.8e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='1.467451345e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.527577506e-07 wvth0=-3.960080134e-07 pvth0=6.183110718e-14 k1=0.90707349 k2=-1.307830464e-01 lk2=-5.033066503e-10 wk2=-3.414267389e-09 pk2=5.330900531e-16 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.585131559e-01 ldsub=1.824357490e-11 wdsub=6.967175620e-11 pdsub=-1.087826933e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.335147271e-19 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749045353e-17 nfactor=6.350352380e+00 lnfactor=-6.051243760e-07 wnfactor=-2.336063788e-06 pnfactor=3.647436557e-13 eta0=1.641773873e-02 leta0=-2.563400019e-09 weta0=-9.789604030e-09 peta0=1.528509615e-15 etab=-0.043998 u0=-1.042515434e-01 lu0=2.081369681e-08 wu0=7.507878410e-08 pu0=-1.172250103e-14 ua=-1.067214387e-09 lua=-1.779247122e-17 wua=-6.809054781e-17 pua=1.063138577e-23 ub=7.948211672e-18 lub=-9.269887297e-25 wub=-3.519397732e-24 pub=5.495046843e-31 uc=3.253499472e-10 luc=-3.877574281e-17 wuc=-1.480842181e-16 puc=2.312127748e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.272164970e+05 lvsat=9.189705032e-03 wvsat=3.365213780e-02 pvsat=-5.254310187e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.700000007e-02 lketa=9.208522833e-18 dwg=0.0 dwb=0.0 pclm=-2.993692922e-01 lpclm=7.474772202e-08 wpclm=2.764238741e-07 ppclm=-4.315971801e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000002e-08 lalpha0=-2.022661738e-24 alpha1=0.85 beta0=1.391835560e+01 lbeta0=-8.622102004e-9 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.708984723e-01 lkt1=3.736038441e-08 wkt1=1.410325905e-07 pkt1=-2.202026454e-14 kt2=-0.028878939 at=5.372048692e+04 lat=1.013628207e-11 ute=2.117734108e-01 lute=-2.385029154e-07 wute=-9.026085853e-07 pute=1.409296941e-13 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.135 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.136 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-7 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-8 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-07 wa0=-7.105427358e-21 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-07 ppclm=8.881784197e-28 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+03 ppscbe1=-1.525878906e-17 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-7 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-6 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.137 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-8 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 wpclm=4.440892099e-22 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-8 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 wuc1=2.067951531e-31 puc1=-8.271806126e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.138 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-06 wdsub=-3.552713679e-21 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-8 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-06 wa0=-7.105427358e-21 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-8 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 pua1=-1.323488980e-35 ub1=-1.486104833e-18 lub1=3.235003467e-24 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.139 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-7 eta0=-1.482776250e-03 leta0=3.918235528e-09 peta0=-6.938893904e-30 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=-1.804112415e-22 petab=1.179611964e-28 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 pua=3.308722450e-36 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-6 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 wketa=5.551115123e-23 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 palpha0=-1.990527426e-32 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-7 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-2 ute=-2.370540520e+00 lute=1.265004727e-6 ua1=-1.560482787e-09 lua1=2.774223792e-15 wua1=-1.654361225e-30 pua1=6.617444900e-36 ub1=9.526220239e-19 lub1=-1.584252469e-24 wub1=-1.540743956e-39 uc1=7.177850760e-11 luc1=-3.002883819e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.140 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.379634364e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.432720057e-8 k1=6.296133047e-01 lk1=-7.362455483e-8 k2=-6.835126213e-02 lk2=2.800349610e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242964e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338157261e-9 nfactor=2.783078619e+00 lnfactor=9.531360947e-8 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=7.355227538e-22 peta0=3.469446952e-28 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.955893720e-02 lu0=-3.867194305e-9 ua=-8.304373631e-10 lua=-2.958561202e-16 ub=1.698955783e-18 lub=9.402944032e-26 uc=2.718870035e-11 luc=1.206923800e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-8.676901760e+02 lvsat=8.227234419e-2 a0=1.024210589e+00 la0=1.715943727e-7 ags=2.291547500e+00 lags=-1.016692010e-6 a1=0.0 a2=0.42385546 b0=2.229104170e-07 lb0=-1.061356743e-13 b1=4.301245670e-09 lb1=-2.047977909e-15 keta=-1.155907111e-01 lketa=5.164999439e-8 dwg=0.0 dwb=0.0 pclm=1.268894400e+00 lpclm=-3.890432980e-7 pdiblc1=6.603681753e-01 lpdiblc1=-2.986974357e-7 pdiblc2=9.120988833e-03 lpdiblc2=-4.320720495e-9 pdiblcb=8.971602892e-02 lpdiblcb=-8.776197741e-08 wpdiblcb=-1.249000903e-22 ppdiblcb=4.770489559e-29 drout=8.432395256e-01 ldrout=7.463925761e-8 pscbe1=1.016674454e+09 lpscbe1=-2.760291061e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680640e-06 lalpha0=-1.505866109e-12 alpha1=0.85 beta0=1.693644131e+01 lbeta0=5.149690275e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693353e-01 lkt1=-3.990136189e-9 kt2=-1.799095058e-02 lkt2=-8.916908084e-9 at=1.122373800e+05 lat=-4.836690427e-2 ute=-8.501885196e-01 lute=-2.190655934e-7 ua1=1.709985088e-09 lua1=-4.181976374e-16 ub1=-7.070069558e-19 lub1=3.577112438e-26 uc1=7.460704526e-11 luc1=-3.278987563e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.141 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.143892664e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.206188842e-8 k1=8.414013971e-02 lk1=1.860948561e-7 k2=1.094279808e-01 lk2=-5.664360154e-08 wk2=5.551115123e-23 pk2=-6.938893904e-29 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425679e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-09 pcdscd=-6.938893904e-30 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663645e-8 nfactor=3.588363944e+00 lnfactor=-2.881117241e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=-4.510281038e-23 petab=2.428612866e-29 u0=1.679523247e-02 lu0=2.210065012e-9 ua=-1.703807103e-09 lua=1.199866543e-16 ub=1.993090003e-18 lub=-4.601845039e-26 uc=1.633443547e-11 luc=1.723734426e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.663999498e+05 lvsat=2.630199184e-3 a0=1.280215623e+00 la0=4.970115984e-8 ags=-8.330949999e-01 lags=4.710627709e-07 wags=1.776356839e-21 pags=4.440892099e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.166340672e-02 lketa=-3.274707227e-08 pketa=-4.163336342e-29 dwg=0.0 dwb=0.0 pclm=6.446949625e-01 lpclm=-9.183947451e-08 wpclm=-3.552713679e-21 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 ppdiblc1=-2.220446049e-28 pdiblc2=-7.515255684e-03 lpdiblc2=3.600394425e-09 wpdiblc2=-5.204170428e-24 ppdiblc2=2.710505431e-30 pdiblcb=-8.674421609e-02 lpdiblcb=-3.742902196e-9 drout=1.449262700e+00 ldrout=-2.139101923e-07 wdrout=-7.105427358e-21 pscbe1=1.163107023e+08 lpscbe1=1.526664890e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183449e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126010e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532692e+03 lat=7.780439669e-03 pat=1.455191523e-23 ute=-1.302351205e+00 lute=-3.774660968e-9 ua1=1.605522255e-09 lua1=-3.684591218e-16 ub1=-1.843635241e-18 lub1=5.769607696e-25 pub1=7.703719778e-46 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=1.550963649e-31 puc1=-3.877409121e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.142 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820499721e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033839681e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217004772e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944755551e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083453410e-16 ags=1.250000000e+00 lags=4.461142566e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566746898e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563738690e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831956891e-18 drout=5.033266588e-01 ldrout=1.889173262e-16 pscbe1=7.914198799e+08 lpscbe1=1.866531372e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.131983396e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135939574e-25 ub1=7.077531681e-19 lub1=3.034217886e-34 uc1=1.471862500e-10 luc1=-4.393156233e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.143 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.4e-07 wmax=5.5e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='-3.172849528e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.717602665e-07 wvth0=1.953292793e-06 pvth0=-3.049793236e-13 k1=0.90707349 k2=-3.003671695e-01 lk2=2.597487998e-08 wk2=8.244312159e-08 pk2=-1.287233923e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.467965476e+00 ldsub=-3.137296038e-07 wdsub=-1.017279868e-06 pdsub=1.588340094e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.335181965e-19 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749000944e-17 nfactor=-2.028325946e+00 lnfactor=7.030889431e-07 wnfactor=1.905910232e-06 pnfactor=-2.975812000e-13 eta0=-1.136608897e-02 leta0=1.774655702e-09 weta0=4.276847823e-09 peta0=-6.677699117e-16 etab=-0.043998 u0=7.908565556e-01 lu0=-1.189449013e-07 wu0=-3.780983345e-07 pu0=5.903476155e-14 ua=-1.477932634e-09 lua=4.633543300e-17 wua=1.398487077e-16 pua=-2.183541783e-23 ub=6.883165008e-18 lub=-7.606966037e-25 wub=-2.980183777e-24 pub=4.653139742e-31 uc=-2.014268080e-10 luc=4.347307263e-17 wuc=1.186133710e-16 puc=-1.851981730e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=9.001357668e+05 lvsat=-1.114908181e-01 wvsat=-3.576629760e-01 pvsat=5.584406642e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.229130883e-01 lketa=1.242706859e-07 wketa=4.029564701e-07 pketa=-6.291601142e-14 dwg=0.0 dwb=0.0 pclm=8.088112420e-03 lpclm=2.674255270e-08 wpclm=1.207637244e-07 ppclm=-1.885556487e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.999997574e-08 lalpha0=3.788690917e-21 walpha0=1.229165593e-20 palpha0=-1.919170088e-27 alpha1=0.85 beta0=1.391835537e+01 lbeta0=-8.622065789e-09 wbeta0=1.174323643e-13 pbeta0=-1.833538477e-20 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.923331776e-01 lkt1=-6.133686455e-09 wkt1=-4.101782025e-15 pkt1=6.404361486e-22 kt2=-0.028878939 at=5.372048954e+04 lat=-3.982814960e-10 wat=-1.324324869e-09 pat=2.067746827e-16 ute=-1.132927112e+00 lute=-2.854675466e-08 wute=-2.218109154e-07 pute=3.463266909e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.144 nmos lmin=2.0e-05 lmax=0.0001 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.145 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.685741570e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.058779873e-7 k1=6.123320250e-01 lk1=-8.854283449e-7 k2=-5.163799463e-02 lk2=3.028991216e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.016862216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.316750651e-7 nfactor=3.665874199e+00 lnfactor=-6.403833805e-6 eta0=0.08 etab=-0.07 u0=2.231223305e-02 lu0=4.094842102e-08 wu0=5.551115123e-23 ua=-1.241809818e-09 lua=3.755336140e-15 ub=1.685065637e-18 lub=-1.765203975e-24 uc=6.330548048e-11 luc=-2.950171746e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.390915283e+00 la0=-5.656299401e-7 ags=3.208651839e-01 lags=4.797232332e-7 a1=0.0 a2=0.42385546 b0=2.422797401e-08 lb0=-1.797800326e-14 b1=5.203866371e-09 lb1=-2.581848400e-14 keta=-2.660376772e-03 lketa=-3.767945174e-8 dwg=0.0 dwb=0.0 pclm=-9.712120000e-03 lpclm=5.311079250e-7 pdiblc1=0.39 pdiblc2=5.516568119e-04 lpdiblc2=8.163660446e-9 pdiblcb=-0.025 drout=0.56 pscbe1=-7.410457490e+07 lpscbe1=5.974953667e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.832161327e-01 lkt1=-6.320184307e-8 kt2=-3.546454717e-02 lkt2=1.187904134e-7 at=1.982637300e+05 lat=-4.647194343e-1 ute=-1.015897703e+00 lute=-1.987671409e-6 ua1=1.029872646e-09 lua1=1.820372413e-15 ub1=-3.826688949e-19 lub1=-3.731564281e-24 uc1=6.931016453e-11 luc1=-7.089890741e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.146 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.119535564e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=5.987799812e-8 k1=4.369481614e-01 lk1=5.134572035e-7 k2=1.478903246e-02 lk2=-2.269318805e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.179982599e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.568029407e-9 nfactor=2.835644582e+00 lnfactor=2.181905348e-7 eta0=0.08 etab=-0.07 u0=2.571876712e-02 lu0=1.377744198e-8 ua=-9.768594712e-10 lua=1.642056141e-15 ub=1.627914685e-18 lub=-1.309360213e-24 uc=9.599342154e-12 luc=1.333502887e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.409463060e+00 la0=-7.135695335e-7 ags=3.609702746e-01 lags=1.598395755e-7 a1=0.0 a2=0.42385546 b0=1.082491466e-08 lb0=8.892662098e-14 b1=5.983139888e-10 lb1=1.091602815e-14 keta=-1.746390476e-02 lketa=8.039550078e-08 pketa=1.110223025e-28 dwg=0.0 dwb=0.0 pclm=-6.945600321e-01 lpclm=5.993548011e-06 wpclm=6.661338148e-22 ppclm=-1.776356839e-27 pdiblc1=0.39 pdiblc2=-1.643357236e-03 lpdiblc2=2.567139102e-08 ppdiblc2=-2.775557562e-29 pdiblcb=-0.025 drout=0.56 pscbe1=6.390114615e+08 lpscbe1=2.870431763e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.862692334e-01 lkt1=-3.884989683e-8 kt2=-9.795153463e-03 lkt2=-8.595216188e-8 at=140000.0 ute=-1.231004634e+00 lute=-2.719492778e-7 ua1=1.515902718e-09 lua1=-2.056269539e-15 wua1=-3.308722450e-30 ub1=-1.027457992e-18 lub1=1.411361252e-24 uc1=-7.120287721e-11 luc1=4.117620565e-16 wuc1=-5.169878828e-32 puc1=2.067951531e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.147 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.356425871e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-3.431280957e-8 k1=5.591506344e-01 lk1=2.756355115e-8 k2=-3.970628007e-02 lk2=-1.025110655e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.564204000e-01 ldsub=-1.178607824e-6 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.372392365e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.493671045e-8 nfactor=2.540960508e+00 lnfactor=1.389894491e-6 eta0=1.585514060e-01 leta0=-3.123310732e-7 etab=-1.386707260e-01 letab=2.730441458e-7 u0=3.009815813e-02 lu0=-3.635612266e-9 ua=-7.055192805e-10 lua=5.631706405e-16 ub=1.674767488e-18 lub=-1.495653328e-24 uc=3.557531560e-11 luc=3.006628558e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.610603794e+00 la0=-1.513332445e-6 ags=3.267882410e-01 lags=2.957519899e-7 a1=0.0 a2=0.42385546 b0=6.450162160e-10 lb0=1.294032816e-13 b1=-1.306345622e-09 lb1=1.848921380e-14 keta=5.179224004e-04 lketa=8.897310460e-9 dwg=0.0 dwb=0.0 pclm=1.116334728e+00 lpclm=-1.206815837e-6 pdiblc1=0.39 pdiblc2=2.474187624e-03 lpdiblc2=9.299472665e-9 pdiblcb=-3.735085000e-02 lpdiblcb=4.910865932e-8 drout=0.56 pscbe1=6.234654264e+08 lpscbe1=3.488563261e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.587107910e-01 lkt1=-1.484260119e-7 kt2=-1.476078455e-02 lkt2=-6.620813734e-8 at=1.702645228e+05 lat=-1.203358588e-1 ute=-8.735426920e-01 lute=-1.693266573e-6 ua1=2.140334125e-09 lua1=-4.539093737e-15 ub1=-1.486104833e-18 lub1=3.235003467e-24 pub1=-6.162975822e-45 uc1=8.417239227e-12 luc1=9.518164525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.148 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.847371124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=6.628333163e-8 k1=5.915575913e-01 lk1=-3.647700292e-8 k2=-4.999948451e-02 lk2=1.008966530e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.26 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-6.481406205e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-6.818528415e-8 nfactor=3.599201184e+00 lnfactor=-7.013330064e-7 eta0=-1.482776250e-03 leta0=3.918235528e-09 peta0=3.469446952e-30 etab=8.137340700e-02 letab=-1.617929870e-07 wetab=2.775557562e-23 petab=-3.122502257e-29 u0=3.085609312e-02 lu0=-5.133394898e-9 ua=2.754445177e-10 lua=-1.375347236e-15 ub=6.147365314e-20 lub=1.692434697e-24 uc=6.175884023e-11 luc=-2.167592006e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=7.666551942e+04 lvsat=6.589387108e-3 a0=4.980764928e-01 la0=6.851728046e-7 ags=-2.786400028e-01 lags=1.492160538e-6 a1=0.0 a2=0.42385546 b0=1.922271293e-08 lb0=9.269122637e-14 b1=1.375707435e-08 lb1=-1.127815269e-14 keta=7.110305558e-02 lketa=-1.305885123e-07 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=1.496432008e-01 lpclm=7.034980908e-7 pdiblc1=4.247813265e-01 lpdiblc1=-6.873263151e-8 pdiblc2=9.606198839e-03 lpdiblc2=-4.794351448e-9 pdiblcb=-2.451476819e-02 lpdiblcb=2.374281595e-8 drout=2.088804448e-01 ldrout=6.938599933e-7 pscbe1=8.645253716e+08 lpscbe1=-1.275109097e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.328986640e-06 lalpha0=1.059008642e-11 walpha0=5.293955920e-28 palpha0=-6.670384460e-33 alpha1=0.85 beta0=1.034200586e+01 lbeta0=6.952034876e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.915711146e-01 lkt1=1.141240567e-7 kt2=-6.889893246e-02 lkt2=4.077620572e-8 at=1.549379515e+05 lat=-9.004846934e-2 ute=-2.370540520e+00 lute=1.265004727e-6 ua1=-1.560482787e-09 lua1=2.774223792e-15 wua1=-1.240770919e-30 pua1=-1.654361225e-36 ub1=9.526220239e-19 lub1=-1.584252469e-24 wub1=7.703719778e-40 pub1=-3.851859889e-46 uc1=7.177850760e-11 luc1=-3.002883819e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.149 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.379634364e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.432720057e-8 k1=6.296133047e-01 lk1=-7.362455483e-8 k2=-6.835126213e-02 lk2=2.800349610e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.120939287e-01 ldsub=4.676284081e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.261242964e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-8.338157261e-9 nfactor=2.783078619e+00 lnfactor=9.531360947e-8 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=-2.636779683e-22 peta0=-4.267419751e-28 etab=-1.641277800e-01 letab=7.784955966e-8 u0=2.955893720e-02 lu0=-3.867194305e-9 ua=-8.304373631e-10 lua=-2.958561202e-16 ub=1.698955783e-18 lub=9.402944032e-26 uc=2.718870035e-11 luc=1.206923800e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-8.676901760e+02 lvsat=8.227234419e-2 a0=1.024210589e+00 la0=1.715943727e-7 ags=2.291547500e+00 lags=-1.016692010e-6 a1=0.0 a2=0.42385546 b0=2.229104170e-07 lb0=-1.061356743e-13 b1=4.301245670e-09 lb1=-2.047977909e-15 keta=-1.155907111e-01 lketa=5.164999439e-8 dwg=0.0 dwb=0.0 pclm=1.268894400e+00 lpclm=-3.890432980e-7 pdiblc1=6.603681753e-01 lpdiblc1=-2.986974357e-7 pdiblc2=9.120988833e-03 lpdiblc2=-4.320720495e-9 pdiblcb=8.971602892e-02 lpdiblcb=-8.776197741e-08 wpdiblcb=-8.413408858e-23 ppdiblcb=1.023486851e-28 drout=8.432395256e-01 ldrout=7.463925761e-8 pscbe1=1.016674454e+09 lpscbe1=-2.760291061e+02 wpscbe1=-1.907348633e-12 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.062680640e-06 lalpha0=-1.505866109e-12 alpha1=0.85 beta0=1.693644131e+01 lbeta0=5.149690275e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.705693353e-01 lkt1=-3.990136189e-9 kt2=-1.799095058e-02 lkt2=-8.916908084e-9 at=1.122373800e+05 lat=-4.836690427e-02 wat=-2.328306437e-16 ute=-8.501885196e-01 lute=-2.190655934e-7 ua1=1.709985088e-09 lua1=-4.181976374e-16 wua1=3.308722450e-30 ub1=-7.070069558e-19 lub1=3.577112438e-26 uc1=7.460704526e-11 luc1=-3.278987563e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.150 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.143892664e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-2.206188842e-8 k1=8.414013971e-02 lk1=1.860948561e-7 k2=1.094279808e-01 lk2=-5.664360154e-08 wk2=-2.775557562e-23 pk2=6.938893904e-30 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.761425679e-01 ldsub=6.388057796e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.121188879e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.500663645e-8 nfactor=3.588363944e+00 lnfactor=-2.881117241e-7 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.860778692e-02 letab=-1.868014223e-08 wetab=2.775557562e-23 petab=5.637851297e-30 u0=1.679523247e-02 lu0=2.210065012e-9 ua=-1.703807103e-09 lua=1.199866543e-16 ub=1.993090003e-18 lub=-4.601845039e-26 uc=1.633443547e-11 luc=1.723734426e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.663999498e+05 lvsat=2.630199184e-3 a0=1.280215623e+00 la0=4.970115984e-8 ags=-8.330949999e-01 lags=4.710627709e-07 wags=4.440892099e-22 pags=4.440892099e-28 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=6.166340672e-02 lketa=-3.274707227e-08 wketa=-2.775557562e-23 pketa=2.081668171e-29 dwg=0.0 dwb=0.0 pclm=6.446949625e-01 lpclm=-9.183947451e-8 pdiblc1=-2.599865133e-01 lpdiblc1=1.395165643e-07 wpdiblc1=-1.110223025e-22 ppdiblc1=2.775557562e-29 pdiblc2=-7.515255684e-03 lpdiblc2=3.600394425e-09 wpdiblc2=2.168404345e-25 ppdiblc2=3.794707604e-31 pdiblcb=-8.674421609e-02 lpdiblcb=-3.742902196e-9 drout=1.449262700e+00 ldrout=-2.139101923e-7 pscbe1=1.163107023e+08 lpscbe1=1.526664890e+2 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=7.408183449e-06 lalpha0=-1.670372435e-12 alpha1=0.85 beta0=2.136300371e+01 lbeta0=-1.592676687e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.133121573e-01 lkt1=1.636126010e-8 kt2=-4.380991832e-02 lkt2=3.376431938e-9 at=-5.685532692e+03 lat=7.780439669e-3 ute=-1.302351205e+00 lute=-3.774660968e-9 ua1=1.605522255e-09 lua1=-3.684591218e-16 ub1=-1.843635241e-18 lub1=5.769607696e-25 uc1=-1.222035414e-10 luc1=6.091872988e-17 wuc1=-1.033975766e-31 puc1=-3.231174268e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.151 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.787058597e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.399258556e-8 k1=9.070734896e-01 lk1=6.820322085e-17 k2=-1.567821040e-01 lk2=3.556082198e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=4.586300001e-01 ldsub=-1.033750863e-17 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999996e-03 lcdscd=7.217039466e-19 cit=0.0 voff='-1.136835598e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280779e-8 nfactor=1.956461452e+00 lnfactor=8.092017789e-8 eta0=2.242428860e-03 leta0=-3.501238375e-10 etab=-4.399800002e-02 letab=2.944755551e-18 u0=2.102562674e-02 lu0=1.253420572e-9 ua=-1.155463028e-09 lua=-4.013681436e-18 ub=1.295395749e-18 lub=1.117553374e-25 uc=1.272578803e-10 luc=-7.846439865e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.600919746e+05 lvsat=4.056659463e-3 a0=1.499999999e+00 la0=2.083488937e-16 ags=1.250000000e+00 lags=4.460964931e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-2.083869161e-01 lketa=2.832102752e-8 dwg=0.0 dwb=0.0 pclm=3.706266759e-01 lpclm=-2.986276845e-8 pdiblc1=3.569721502e-01 lpdiblc1=-3.566924534e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563599912e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831734847e-18 drout=5.033266588e-01 ldrout=1.889155499e-16 pscbe1=7.914198799e+08 lpscbe1=1.866149902e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=2.863680696e-09 lalpha0=4.236956351e-15 alpha1=0.85 beta0=1.533904646e+01 lbeta0=-2.304430895e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.618011205e-01 lkt1=4.712760272e-9 kt2=-2.887893901e-02 lkt2=1.131983396e-18 at=-2.704237011e+04 lat=1.260998945e-2 ute=-1.326367013e+00 lute=1.656177765e-9 ua1=-2.384733737e-11 lua1=2.135940608e-25 ub1=7.077531681e-19 lub1=3.034187072e-34 uc1=1.471862500e-10 luc1=-4.393363028e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.152 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=5.2e-07 wmax=5.4e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='2.525953477e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.692500534e-08 wvth0=2.533061593e-07 pvth0=-3.955021049e-14 k1=0.90707349 k2=-1.842726492e-01 lk2=7.848345977e-09 wk2=2.482750091e-08 pk2=-3.876466683e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.467965459e+00 ldsub=-3.137296012e-07 wdsub=-1.017279859e-06 pdsub=1.588340081e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000001e-03 lcdscd=-1.335112576e-19 cit=0.0 voff='-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.749089762e-17 nfactor=-2.028325776e+00 lnfactor=7.030889166e-07 wnfactor=1.905910148e-06 pnfactor=-2.975811868e-13 eta0=-1.136614629e-02 leta0=1.774664653e-09 weta0=4.276876273e-09 peta0=-6.677743538e-16 etab=-0.043998 u0=6.262738395e-02 lu0=-5.242111391e-09 wu0=-1.669130470e-08 pu0=2.606113551e-15 ua=-1.477932599e-09 lua=4.633542753e-17 wua=1.398486904e-16 pua=-2.183541512e-23 ub=6.883164335e-18 lub=-7.606964985e-25 wub=-2.980183442e-24 pub=4.653139219e-31 uc=-2.014268208e-10 luc=4.347307463e-17 wuc=1.186133774e-16 puc=-1.851981829e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.736637301e+05 lvsat=-1.367598016e-02 wvsat=-4.675618067e-02 pvsat=7.300323024e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-8.229130756e-01 lketa=1.242706840e-07 wketa=4.029564638e-07 pketa=-6.291601043e-14 dwg=0.0 dwb=0.0 pclm=8.088139166e-03 lpclm=2.674254852e-08 wpclm=1.207637111e-07 ppclm=-1.885556280e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.000000006e-08 lalpha0=-9.450452472e-24 walpha0=2.191735868e-22 palpha0=-3.422087222e-29 alpha1=0.85 beta0=1.391835560e+01 lbeta0=-8.622102722e-09 wbeta0=3.967670636e-17 pbeta0=-6.210143511e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.923331857e-01 lkt1=-6.133685191e-09 wkt1=-8.154366071e-17 pkt1=1.273181560e-23 kt2=-0.028878939 at=5.372048692e+04 lat=1.022242941e-11 wat=-2.588424832e-11 pat=4.041474313e-18 ute=-1.132927148e+00 lute=-2.854674899e-08 wute=-2.218108973e-07 pute=3.463266627e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.153 nmos lmin=2.0e-05 lmax=0.0001 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.154 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.440467258e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=8.958412891e-07 wvth0=1.168197400e-08 pvth0=-2.333607013e-13 k1=8.217577412e-01 lk1=-5.068944934e-06 wk1=-9.974569897e-08 pk1=1.992533648e-12 k2=-1.408123644e-01 lk2=2.084258460e-06 wk2=4.247214719e-08 pk2=-8.484293884e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.014047019e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.372987414e-07 wvoff=-1.340827786e-10 pvoff=2.678455820e-15 nfactor=4.247871716e+00 lnfactor=-1.802989535e-05 wnfactor=-2.771949411e-07 pnfactor=5.537283843e-12 eta0=0.08 etab=-0.07 u0=1.906185070e-02 lu0=1.058785009e-07 wu0=1.548098606e-09 pu0=-3.092502829e-14 ua=-1.616986101e-09 lua=1.124990859e-14 wua=1.786897104e-16 pua=-3.569529956e-21 ub=1.862903844e-18 lub=-5.317724193e-24 wub=-8.470113711e-26 pub=1.692001434e-30 uc=6.326296240e-11 luc=-2.941678276e-16 wuc=2.025059733e-20 puc=-4.045286864e-25 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.060774878e+00 la0=6.029299683e-06 wa0=1.572399322e-07 pa0=-3.141046271e-12 ags=3.186892585e-01 lags=5.231898148e-07 wags=1.036354099e-09 pags=-2.070235042e-14 a1=0.0 a2=0.42385546 b0=6.783401913e-08 lb0=-8.890582910e-13 wb0=-2.076877438e-14 pb0=4.148798616e-19 b1=8.875177735e-09 lb1=-9.915709911e-14 wb1=-1.748579519e-15 pb1=3.492986228e-20 keta=-5.263483841e-03 lketa=1.432056911e-08 wketa=1.239813041e-09 pketa=-2.476667393e-14 dwg=0.0 dwb=0.0 pclm=5.695623324e-02 lpclm=-8.006681662e-07 wpclm=-3.175293662e-08 ppclm=6.343009803e-13 pdiblc1=0.39 pdiblc2=3.210332764e-03 lpdiblc2=-4.494641196e-08 wpdiblc2=-1.266279500e-09 ppdiblc2=2.529537151e-14 pdiblcb=-0.025 drout=0.56 pscbe1=-1.041850928e+08 lpscbe1=6.575846183e+03 wpscbe1=1.432680922e+01 ppscbe1=-2.861942893e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.009236635e-01 lkt1=2.905262004e-07 wkt1=8.433778183e-09 pkt1=-1.684743000e-13 kt2=-6.178975046e-02 lkt2=6.446662545e-07 wkt2=1.253822047e-08 pkt2=-2.504651974e-13 at=2.357796851e+05 lat=-1.214143255e+00 wat=-1.786817412e-02 pat=3.569370762e-7 ute=-6.094748567e-01 lute=-1.010642947e-05 wute=-1.935718863e-07 pute=3.866818326e-12 ua1=1.606117716e-09 lua1=-9.690777475e-15 wua1=-2.744551544e-16 pua1=5.482553491e-21 ub1=-8.876086396e-19 lub1=6.355180732e-24 wub1=2.404937115e-25 pub1=-4.804135088e-30 uc1=1.677082470e-10 luc1=-2.674602552e-15 wuc1=-4.686523553e-17 puc1=9.361863187e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.155 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.204799510e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=2.861994897e-07 wvth0=-4.060968279e-09 pvth0=-1.077928527e-13 k1=-2.040130716e-01 lk1=3.112742574e-06 wk1=3.052782980e-07 pk1=-1.237992835e-12 k2=2.880568093e-01 lk2=-1.336460396e-06 wk2=-1.301525233e-07 pk2=5.284484603e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-8.790875386e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.449442585e-07 wvoff=-1.433109012e-08 pvoff=1.159157171e-13 nfactor=1.543659763e+00 lnfactor=3.539266966e-06 wnfactor=6.153491137e-07 pnfactor=-1.581768925e-12 eta0=0.08 etab=-0.07 u0=3.156833316e-02 lu0=6.125095903e-09 wu0=-2.786043012e-09 pu0=3.644674696e-15 ua=-1.865050936e-11 lua=-1.498633460e-15 wua=-4.563776808e-16 pua=1.495853925e-21 ub=9.153859060e-19 lub=2.239807743e-24 wub=3.393646320e-25 pub=-1.690404813e-30 uc=-7.681406779e-11 luc=8.231056157e-16 wuc=4.115715172e-17 puc=-3.285180466e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=2.175462013e+00 la0=-2.861596503e-06 wa0=-3.648315134e-07 pa0=1.023066581e-12 ags=1.893441793e-01 lags=1.554863758e-06 wags=8.174241992e-08 pags=-6.644249075e-13 a1=0.0 a2=0.42385546 b0=-2.289842658e-07 lb0=1.478404717e-12 wb0=1.142167961e-13 pb0=-6.617834064e-19 b1=-1.292107121e-09 lb1=-1.806145234e-14 wb1=9.003735472e-16 pb1=1.380145237e-20 keta=-1.077482467e-02 lketa=5.827977310e-08 wketa=-3.185888443e-09 pketa=1.053332301e-14 dwg=0.0 dwb=0.0 pclm=-2.008746810e+00 lpclm=1.567566024e-05 wpclm=6.259235070e-07 ppclm=-4.611415778e-12 pdiblc1=0.39 pdiblc2=-3.884875667e-03 lpdiblc2=1.164593544e-08 wpdiblc2=1.067594881e-09 ppdiblc2=6.680072035e-15 pdiblcb=-0.025 drout=0.56 pscbe1=1.061386927e+09 lpscbe1=-2.720914767e+03 wpscbe1=-2.011698316e+02 ppscbe1=1.432636225e-3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.995756302e-01 lkt1=2.797741037e-07 wkt1=6.337597304e-09 pkt1=-1.517548762e-13 kt2=2.322492653e-02 lkt2=-3.342237117e-08 wkt2=-1.572686974e-08 pkt2=-2.501899378e-14 at=2.745213476e+04 lat=4.475056187e-01 wat=5.360452235e-02 pat=-2.131388711e-7 ute=-2.827302572e+00 lute=7.583266016e-06 wute=7.602879747e-07 pute=-3.741297650e-12 ua1=-1.784648604e-09 lua1=1.735443584e-14 wua1=1.571993185e-15 pua1=-9.244969580e-21 ub1=1.459670687e-18 lub1=-1.236703841e-23 wub1=-1.184574622e-24 pub1=6.562403748e-30 uc1=-2.939811106e-10 luc1=1.007894554e-15 wuc1=1.061052626e-16 puc1=-2.839271782e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.156 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.381992291e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.818683698e-07 wvth0=-4.884588258e-08 pvth0=7.027805733e-14 k1=6.989797175e-01 lk1=-4.776795624e-07 wk1=-6.659807534e-08 pk1=2.406382006e-13 k2=-1.061923299e-01 lk2=2.311277994e-07 wk2=3.166610877e-08 pk2=-1.149644281e-13 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.971797010e+00 ldsub=-5.613496914e-06 wdsub=-5.312338023e-07 pdsub=2.112257846e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-2.337651669e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=3.350006763e-07 wvoff=4.597356318e-08 pvoff=-1.238637858e-13 nfactor=1.568996789e+00 lnfactor=3.438523505e-06 wnfactor=4.629288240e-07 pnfactor=-9.757251240e-13 eta0=4.541262075e-01 leta0=-1.487576682e-06 weta0=-1.407769576e-07 peta0=5.597483292e-13 etab=-3.970663072e-01 letab=1.300460118e-06 wetab=1.230691642e-07 petab=-4.893397343e-13 u0=3.560475970e-02 lu0=-9.924284997e-09 wu0=-2.622695211e-09 pu0=2.995181625e-15 ua=-1.503415702e-09 lua=4.404994874e-15 wua=3.800237035e-16 pua=-1.829791730e-21 ub=3.565806593e-18 lub=-8.298625364e-24 wub=-9.006678870e-25 pub=3.240133127e-30 uc=1.888221299e-10 luc=-2.331000331e-16 wuc=-7.298869923e-17 puc=1.253413806e-22 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.328186982e+05 lvsat=-1.005241527e+00 wvsat=-1.204129952e-01 pvsat=4.787784451e-7 a0=4.495430831e+00 la0=-1.208610804e-05 wa0=-1.373991191e-06 pa0=5.035622705e-12 ags=-9.049205322e-02 lags=2.667530676e-06 wags=1.987430931e-07 pags=-1.129635496e-12 a1=0.0 a2=0.42385546 b0=-9.209822745e-08 lb0=9.341272118e-13 wb0=4.417193758e-14 pb0=-3.832755229e-19 b1=-1.914328479e-08 lb1=5.291725781e-14 wb1=8.495413059e-15 pb1=-1.639745766e-20 keta=5.073748949e-02 lketa=-1.863015537e-07 wketa=-2.391867585e-08 pketa=9.296970541e-14 dwg=0.0 dwb=0.0 pclm=8.147361128e+00 lpclm=-2.470640615e-05 wpclm=-3.348751316e-06 ppclm=1.119243187e-11 pdiblc1=0.39 pdiblc2=1.418717630e-02 lpdiblc2=-6.021100098e-08 wpdiblc2=-5.578685672e-09 ppdiblc2=3.310658741e-14 pdiblcb=-8.382487540e-02 lpdiblcb=2.338957048e-07 wpdiblcb=2.213474176e-08 ppdiblcb=-8.801074358e-14 drout=0.56 pscbe1=-4.080239783e+07 lpscbe1=1.661539887e+03 wpscbe1=3.163788079e+02 ppscbe1=-6.252075519e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-8.194415328e-02 lkt1=-5.855582466e-07 wkt1=-8.419076773e-08 pkt1=2.081982150e-13 kt2=1.434144464e-01 lkt2=-5.113122478e-07 wkt2=-7.533601533e-08 pkt2=2.119950759e-13 at=2.841444747e+05 lat=-5.731380349e-01 wat=-5.423897122e-02 pat=2.156615261e-7 ute=1.909014365e+00 lute=-1.124897427e-05 wute=-1.325281840e-06 pute=4.551211572e-12 ua1=1.141786848e-08 lua1=-3.514056761e-14 wua1=-4.418722615e-15 pua1=1.457493118e-20 ub1=-7.308256149e-18 lub1=2.249543113e-23 wub1=2.772985873e-24 pub1=-9.173395008e-30 uc1=-1.786418358e-10 luc1=5.492899110e-16 wuc1=8.909287036e-17 puc1=-2.162835930e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.157 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.504369097e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.891755091e-07 wvth0=1.633656913e-08 pvth0=-5.853133206e-14 k1=4.780953274e-01 lk1=-4.118196720e-08 wk1=5.404003399e-08 pk1=2.240889795e-15 k2=2.993537022e-03 lk2=1.536167717e-08 wk2=-2.523962228e-08 pk2=-2.510964359e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-1.970753219e+00 ldsub=2.177518524e-06 wdsub=1.062467605e-06 pdsub=-1.037112878e-12 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='5.996276874e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.454456715e-07 wvoff=-5.942895852e-08 pvoff=8.442593182e-14 nfactor=5.245328609e+00 lnfactor=-3.826408152e-06 wnfactor=-7.840208619e-07 pnfactor=1.488417041e-12 eta0=-5.926323793e-01 leta0=5.809606445e-07 weta0=2.815539152e-07 peta0=-2.748349126e-13 etab=9.069281548e-01 letab=-1.276410282e-06 wetab=-3.931968664e-07 petab=5.308721543e-13 u0=2.745634634e-02 lu0=6.178087996e-09 wu0=1.619238199e-09 pu0=-5.387455696e-15 ua=2.205141162e-09 lua=-2.923617852e-15 wua=-9.190797770e-16 pua=7.374134259e-22 ub=-3.228910931e-18 lub=5.128660546e-24 wub=1.567150951e-24 pub=-1.636612520e-30 uc=1.124040642e-10 luc=-8.208754232e-17 wuc=-2.412140857e-17 puc=2.877296827e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-8.890861700e+04 lvsat=-1.718509976e-01 wvsat=7.885998084e-02 pvsat=8.498794329e-8 a0=-3.271981319e+00 la0=3.263354737e-06 wa0=1.795610675e-06 pa0=-1.227941647e-12 ags=-2.579801431e+00 lags=7.586744551e-06 wags=1.096001767e-06 pags=-2.902740663e-12 a1=0.0 a2=0.42385546 b0=-6.285731418e-07 lb0=1.994274603e-12 wb0=3.085335053e-13 pb0=-9.056899339e-19 b1=2.303330930e-08 lb1=-3.042942811e-14 wb1=-4.418103732e-15 pb1=9.121407760e-21 keta=2.707199972e-01 lketa=-6.210169064e-07 wketa=-9.507395617e-08 pketa=2.335822164e-13 dwg=0.0 dwb=0.0 pclm=-8.849413375e+00 lpclm=8.881531828e-06 wpclm=4.286088664e-06 ppclm=-3.895050265e-12 pdiblc1=1.288078434e+00 lpdiblc1=-1.774725125e-06 wpdiblc1=-4.111728731e-07 ppdiblc1=8.125335167e-13 pdiblc2=-3.255705279e-02 lpdiblc2=3.216195292e-08 wpdiblc2=2.008159781e-08 ppdiblc2=-1.760162256e-14 pdiblcb=-2.268892823e-02 lpdiblcb=1.130827587e-07 wpdiblcb=-8.696147089e-10 ppdiblcb=-4.255100660e-14 drout=-7.662332490e-01 ldrout=2.620817268e-06 wdrout=4.644291003e-07 pdrout=-9.177750646e-13 pscbe1=1.107322730e+09 lpscbe1=-6.073115110e+02 wpscbe1=-1.156400116e+02 ppscbe1=2.285203900e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-2.549388875e-05 lalpha0=5.043867542e-11 walpha0=9.604179906e-12 palpha0=-1.897916566e-17 alpha1=0.85 beta0=-2.895572869e+00 lbeta0=3.311129075e-05 wbeta0=6.304820470e-06 pbeta0=-1.245918270e-11 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-5.576948819e-01 lkt1=3.545898952e-07 wkt1=7.912176010e-08 pkt1=-1.145295505e-13 kt2=-1.989770592e-01 lkt2=1.652999325e-07 wkt2=6.195387037e-08 pkt2=-5.930840963e-14 at=1.744165334e+05 lat=-3.563006999e-01 wat=-9.277297948e-03 pat=1.268111449e-7 ute=-5.121844387e+00 lute=2.644958824e-06 wute=1.310396508e-06 pute=-6.572472969e-13 ua1=-1.047559365e-08 lua1=8.123891057e-15 wua1=4.246106832e-15 pua1=-2.547950225e-21 ub1=6.164193080e-18 lub1=-4.127960800e-24 wub1=-2.482177486e-24 pub1=1.211522491e-30 uc1=1.802776565e-10 luc1=-1.599838187e-16 wuc1=-5.167619164e-17 puc1=6.189521805e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.158 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.213093526e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.238076616e-08 wvth0=-3.969615964e-08 pvth0=-3.835768323e-15 k1=7.588584447e-01 lk1=-3.152449535e-07 wk1=-6.155713377e-08 pk1=1.150794467e-13 k2=-8.527197030e-02 lk2=1.015208164e-07 wk2=8.059028726e-09 pk2=-3.501497636e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.938772269e-01 ldsub=6.454481925e-08 wdsub=8.676287172e-09 pdsub=-8.469236255e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.993374745e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=7.666630677e-09 wvoff=3.487011889e-08 pvoff=-7.622792408e-15 nfactor=1.595825171e+00 lnfactor=-2.639964645e-07 wnfactor=5.654674471e-07 pnfactor=1.711329207e-13 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=4.336808690e-23 peta0=-1.214306433e-29 etab=-7.805351919e-01 letab=3.707834397e-07 wetab=2.935837549e-07 petab=-1.395191343e-13 u0=5.295665158e-02 lu0=-1.871367796e-08 wu0=-1.114391020e-08 pu0=7.071112928e-15 ua=8.824727399e-10 lua=-1.632513590e-15 wua=-8.158282496e-16 pua=6.366258930e-22 ub=9.981098225e-19 lub=1.002513415e-24 wub=3.338003158e-25 pub=-4.326945643e-31 uc=-1.672334365e-10 luc=1.908766891e-16 wuc=9.259976419e-17 puc=-8.516277042e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-6.554386270e+05 lvsat=3.811593403e-01 wvsat=3.117603549e-01 pvsat=-1.423544963e-7 a0=-7.660993235e-01 la0=8.172731101e-07 wa0=8.526923856e-07 pa0=-3.075251604e-13 ags=9.498328034e+00 lags=-4.203152431e-06 wags=-3.432459846e-06 pags=1.517653742e-12 a1=0.0 a2=0.42385546 b0=2.761403462e-06 lb0=-1.314803599e-12 wb0=-1.209038544e-12 pb0=5.756667763e-19 b1=-1.589157142e-08 lb1=7.566549250e-15 wb1=9.617475310e-15 pb1=-4.579226224e-21 keta=-6.875240046e-01 lketa=3.143595604e-07 wketa=2.724015329e-07 pketa=-1.251238375e-13 dwg=0.0 dwb=0.0 pclm=6.631978465e-01 lpclm=-4.040704387e-07 wpclm=2.884823660e-07 ppclm=7.157156668e-15 pdiblc1=6.058912244e-01 lpdiblc1=-1.108817631e-06 wpdiblc1=2.594639114e-08 ppdiblc1=3.858456666e-13 pdiblc2=5.300944978e-03 lpdiblc2=-4.792601592e-09 wpdiblc2=1.819418127e-09 ppdiblc2=2.247484731e-16 pdiblcb=5.213717968e-01 lpdiblcb=-4.179945013e-07 wpdiblcb=-2.055898725e-07 ppdiblcb=1.572838069e-13 drout=2.793467272e+00 ldrout=-8.539345596e-07 wdrout=-9.288583713e-07 pdrout=4.422629948e-13 pscbe1=1.831981422e+09 lpscbe1=-1.314676947e+03 wpscbe1=-3.883160333e+02 ppscbe1=4.946892711e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.556783204e-05 lalpha0=-9.165868466e-12 walpha0=-1.357649052e-11 palpha0=3.648321242e-18 alpha1=0.85 beta0=3.474735315e+01 lbeta0=-3.633324486e-06 wbeta0=-8.483016712e-06 pbeta0=1.975757531e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.102434031e-01 lkt1=1.542999846e-08 wkt1=-2.873215566e-08 pkt1=-9.249460571e-15 kt2=-7.005837389e-02 lkt2=3.945776265e-08 wkt2=2.479877651e-08 pkt2=-2.303998493e-14 at=-4.204198185e+05 lat=2.243404773e-01 wat=2.536950358e-01 pat=-1.298856171e-7 ute=-4.085857808e+00 lute=1.633695028e-06 wute=1.541091040e-06 pute=-8.824365344e-13 ua1=-6.618614713e-09 lua1=4.358955067e-15 wua1=3.966762170e-15 pua1=-2.275271845e-21 ub1=6.834047212e-18 lub1=-4.781829534e-24 wub1=-3.591668361e-24 pub1=2.294536477e-30 uc1=3.869173814e-10 luc1=-3.616922933e-16 wuc1=-1.487477915e-16 puc1=1.566503013e-22 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.159 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='8.053394933e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-6.524260893e-08 wvth0=-9.094615596e-08 pvth0=2.056619992e-14 k1=-6.361883992e-01 lk1=3.489870706e-07 wk1=3.430795172e-07 pk1=-7.758262970e-14 k2=3.712710289e-01 lk2=-1.158557411e-07 wk2=-1.247111306e-07 pk2=2.820167624e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.125759715e-01 ldsub=5.564167380e-08 wdsub=-1.735257434e-08 pdsub=3.924041752e-15 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413313e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-1.875374552e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=2.048216691e-09 wvoff=3.592050608e-08 pvoff=-8.122919563e-15 nfactor=-1.100527839e-01 lnfactor=5.482334412e-07 wnfactor=1.761489316e-06 pnfactor=-3.983361480e-13 eta0=9.325986798e-01 leta0=-2.107371650e-7 etab=3.636826934e-02 letab=-1.817370668e-08 wetab=1.066641912e-09 petab=-2.412061354e-16 u0=1.971274378e-03 lu0=5.562295598e-09 wu0=7.060384407e-09 pu0=-1.596607088e-15 ua=-3.788124322e-09 lua=5.913258131e-16 wua=9.927227740e-16 pua=-2.244903572e-22 ub=4.292233931e-18 lub=-5.659376619e-25 wub=-1.095040869e-24 pub=2.476281619e-31 uc=3.612787256e-10 luc=-6.076697773e-17 wuc=-1.642907564e-16 puc=3.715205449e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.152887838e+05 lvsat=1.418827382e-02 wvsat=2.434332837e-02 pvsat=-5.504902904e-9 a0=4.532065711e-01 la0=2.367176788e-07 wa0=3.938895252e-07 pa0=-8.907260166e-14 ags=1.466939411e-01 lags=2.494972189e-07 wags=-4.666558364e-07 pags=1.055276842e-13 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.322954847e-02 lketa=-2.405579330e-08 wketa=1.830535488e-08 pketa=-4.139499730e-15 dwg=0.0 dwb=0.0 pclm=-5.689893378e-01 lpclm=1.826182384e-07 wpclm=5.780559859e-07 ppclm=-1.307192684e-13 pdiblc1=-3.604221043e+00 lpdiblc1=8.957683838e-07 wpdiblc1=1.592798710e-06 ppdiblc1=-3.601891291e-13 pdiblc2=-1.667822168e-02 lpdiblc2=5.672470903e-09 wpdiblc2=4.364155770e-09 ppdiblc2=-9.868927293e-16 pdiblcb=-5.855669086e-01 lpdiblcb=1.090588662e-07 wpdiblcb=2.375802696e-07 ppdiblcb=-5.372545186e-14 drout=1.449261983e+00 ldrout=-2.139100303e-07 wdrout=3.413254115e-13 pdrout=-7.718596329e-20 pscbe1=-2.485492668e+09 lpscbe1=7.410278960e+02 wpscbe1=1.239192113e+03 ppscbe1=-2.802259477e-4 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.105748909e-05 lalpha0=-7.018331815e-12 walpha0=-1.126373859e-11 palpha0=2.547136789e-18 alpha1=0.85 beta0=3.869149493e+01 lbeta0=-5.511272379e-06 wbeta0=-8.253248456e-06 pbeta0=1.866356593e-12 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.207382264e-01 lkt1=-2.718663834e-08 wkt1=-9.171949695e-08 pkt1=2.074108016e-14 kt2=5.052406597e-02 lkt2=-1.795587793e-08 wkt2=-4.492957870e-08 pkt2=1.016019521e-14 at=7.067492197e+04 lat=-9.487408107e-03 wat=-3.636911007e-02 pat=8.224365075e-9 ute=-5.378324727e-02 lute=-2.861208247e-07 wute=-5.946704441e-07 pute=1.344763955e-13 ua1=4.851948294e-09 lua1=-1.102592921e-15 wua1=-1.546214287e-15 pua1=3.496547140e-22 ub1=-6.751768404e-18 lub1=1.686866370e-24 wub1=2.337655479e-24 pub1=-5.286280594e-31 uc1=-8.430044351e-10 luc1=2.239177608e-16 wuc1=3.433044912e-16 puc1=-7.763350443e-23 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.25e-6 sbref=1.24e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.160 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='2.061653274e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=7.025224025e-08 wvth0=1.774343498e-07 pvth0=-4.012429413e-14 k1=9.070734896e-01 lk1=6.820277676e-17 k2=-2.358598238e-01 lk2=2.143840146e-08 wk2=3.766329457e-08 pk2=-8.517026781e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.844318224e+00 ldsub=-3.133539921e-07 wdsub=-6.599783585e-07 pdsub=1.492448661e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999994e-03 lcdscd=1.107712880e-18 wcdscd=8.130007084e-19 pcdscd=-1.838485961e-25 cit=0.0 voff='-1.136835596e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.465280784e-08 wvoff=-1.065039168e-16 pvoff=2.408440114e-23 nfactor=-9.894057697e+00 lnfactor=2.760749176e-06 wnfactor=5.644188962e-06 pnfactor=-1.276354315e-12 eta0=2.242427202e-03 leta0=-3.501234117e-10 weta0=8.967860577e-16 peta0=-2.027956119e-22 etab=-4.399800002e-02 letab=2.944838817e-18 u0=-1.851454145e-02 lu0=1.019487605e-08 wu0=1.883227039e-08 pu0=-4.258654297e-15 ua=-1.020055485e-09 lua=-3.463420164e-17 wua=-6.449217553e-17 pua=1.458400261e-23 ub=6.725316299e-19 lub=2.526073378e-25 wub=2.966589683e-25 pub=-6.708527246e-32 uc=2.485790391e-10 luc=-3.528152142e-17 wuc=-5.778308413e-17 puc=1.306683551e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.408925022e+05 lvsat=8.398351336e-03 wvsat=9.144363076e-03 pvsat=-2.067869689e-9 a0=1.499999999e+00 la0=2.083475614e-16 ags=1.250000000e+00 lags=4.460964931e-17 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-5.556566672e-01 lketa=1.068512200e-07 wketa=1.653983316e-07 pketa=-3.740251712e-14 dwg=0.0 dwb=0.0 pclm=3.856047518e-01 lpclm=-3.324985063e-08 wpclm=-7.133787964e-09 ppclm=1.613206275e-15 pdiblc1=3.569721502e-01 lpdiblc1=-3.566869022e-17 pdiblc2=8.406112094e-03 lpdiblc2=9.563565218e-19 pdiblcb=-1.032957700e-01 lpdiblcb=2.831734847e-18 drout=5.033266588e-01 ldrout=1.889159940e-16 pscbe1=7.914198799e+08 lpscbe1=1.866316795e-8 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.841529940e-07 lalpha0=-3.675908380e-14 walpha0=-8.634483671e-14 palpha0=1.952567599e-20 alpha1=0.85 beta0=1.984497675e+01 lbeta0=-1.249396142e-06 wbeta0=-2.146093491e-06 pbeta0=4.853089976e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.723592454e-01 lkt1=-1.551326758e-08 wkt1=-4.259955513e-08 pkt1=9.633292999e-15 kt2=-2.887893901e-02 lkt2=1.132025029e-18 at=-1.109726076e+05 lat=3.158963765e-02 wat=3.997446138e-02 pat=-9.039664800e-9 ute=-1.018204252e+00 lute=-6.803051626e-08 wute=-1.467723759e-07 pute=3.319051800e-14 ua1=-2.384733737e-11 lua1=2.135939962e-25 ub1=7.077531681e-19 lub1=3.034206331e-34 uc1=1.471862500e-10 luc1=-4.393363028e-27 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.161 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=4.2e-07 wmax=5.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='1.442666050e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-1.228100366e-07 wvth0=-3.135030950e-07 pvth0=3.652871475e-14 k1=0.90707349 k2=-5.135550875e-03 lk2=-1.458596362e-08 wk2=-6.049227457e-08 pk2=6.808591163e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-7.653070645e-01 ldsub=9.410246186e-08 wdsub=5.226696447e-07 pdsub=-3.540906255e-14 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.052000005e-03 lcdscd=-6.359062582e-19 wcdscd=-1.896999918e-18 pcdscd=2.392799500e-25 cit=0.0 voff='-2.075300007e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=8.330447443e-17 wvoff=2.485092132e-16 pvoff=-3.134598137e-23 nfactor=2.562288561e+01 lnfactor=-2.784724284e-06 wnfactor=-1.126386412e-05 pnfactor=1.363601460e-12 eta0=-1.136614502e-02 leta0=1.774664763e-09 weta0=4.276876208e-09 peta0=-6.677744065e-16 etab=-0.043998 u0=1.518526513e-01 lu0=-1.640557596e-08 wu0=-5.918769347e-08 pu0=7.923070781e-15 ua=-1.793883530e-09 lua=8.618821411e-17 wua=2.903304318e-16 pua=-4.081658001e-23 ub=8.336513898e-18 lub=-9.440161977e-25 wub=-3.672387679e-24 pub=5.526257949e-31 uc=-4.845095256e-10 luc=7.917999472e-17 wuc=2.534405742e-16 puc=-3.552638160e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.951236289e+05 lvsat=-1.568267986e-02 wvsat=-5.697714417e-02 pvsat=8.256077967e-9 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.261698858e-02 lketa=2.206317671e-08 wketa=1.702702291e-08 pketa=-1.423641446e-14 dwg=0.0 dwb=0.0 pclm=-2.686070209e-02 lpclm=3.115085549e-08 wpclm=1.374092151e-07 ppclm=-2.095516005e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-3.930083952e-07 lalpha0=5.335658687e-14 walpha0=2.014712848e-13 palpha0=-2.541278195e-20 alpha1=0.85 beta0=3.404518278e+00 lbeta0=1.317551282e-06 wbeta0=5.007551470e-06 pbeta0=-6.316325119e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-4.010308949e-01 lkt1=2.019060909e-08 wkt1=9.939896227e-08 pkt1=-1.253778751e-14 kt2=-0.028878939 at=2.495577075e+05 lat=-2.470212364e-02 wat=-9.327374313e-02 pat=1.176517686e-8 ute=-1.851973592e+00 lute=6.215089330e-08 wute=1.206579809e-07 pute=-8.564988193e-15 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.162 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.163 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.750925212e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.756662574e-07 wvth0=-4.440892099e-22 k1=5.566754387e-01 lk1=2.263751931e-7 k2=-2.793918103e-02 lk2=-1.705116018e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017610378e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.301805274e-7 nfactor=3.511203629e+00 lnfactor=-3.314113452e-6 eta0=0.08 etab=-0.07 u0=2.317604858e-02 lu0=2.369272453e-8 ua=-1.142103671e-09 lua=1.763592594e-15 ub=1.637803688e-18 lub=-8.210928520e-25 wub=-1.540743956e-39 uc=6.331678001e-11 luc=-2.952428955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.478652779e+00 la0=-2.318286092e-6 ags=3.214434537e-01 lags=4.681716359e-7 a1=0.0 a2=0.42385546 b0=1.263931308e-08 lb0=2.135186635e-13 b1=4.228185535e-09 lb1=-6.328150926e-15 keta=-1.968579909e-03 lketa=-5.149887994e-8 dwg=0.0 dwb=0.0 pclm=-2.742977677e-02 lpclm=8.850382462e-7 pdiblc1=0.39 pdiblc2=-1.549079328e-04 lpdiblc2=2.227809388e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.611043278e+07 lpscbe1=5.815261596e+03 ppscbe1=-1.907348633e-18 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.785102125e-01 lkt1=-1.572079458e-7 kt2=-2.846841042e-02 lkt2=-2.096536584e-8 at=1.882935600e+05 lat=-2.655539625e-1 ute=-1.123907878e+00 lute=1.699545360e-7 ua1=8.767308350e-10 lua1=4.879554061e-15 ub1=-2.484770535e-19 lub1=-6.412198755e-24 uc1=4.316007430e-11 luc1=-1.866113153e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.164 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.096875978e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-2.687778576e-10 k1=6.072888189e-01 lk1=-1.773240112e-7 k2=-5.783410041e-02 lk2=6.793434087e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.259947907e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.311118168e-8 nfactor=3.179000049e+00 lnfactor=-6.644125212e-7 eta0=0.08 etab=-0.07 u0=2.416419740e-02 lu0=1.581111515e-8 ua=-1.231511291e-09 lua=2.476719931e-15 ub=1.817275000e-18 lub=-2.252580446e-24 uc=3.256440823e-11 luc=-4.995779590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.205892612e+00 la0=-1.427139067e-7 ags=4.065813044e-01 lags=-2.108994399e-7 a1=0.0 a2=0.42385546 b0=7.455615358e-08 lb0=-2.803384769e-13 b1=1.100708765e-09 lb1=1.861702913e-14 keta=-1.924158216e-02 lketa=8.627293517e-08 pketa=5.551115123e-29 dwg=0.0 dwb=0.0 pclm=-3.453042139e-01 lpclm=3.420447988e-06 ppclm=4.440892099e-28 pdiblc1=0.39 pdiblc2=-1.047655494e-03 lpdiblc2=2.939876984e-8 pdiblcb=-0.025 drout=0.56 pscbe1=5.267617483e+08 lpscbe1=1.086432449e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.827329503e-01 lkt1=-1.235268148e-7 kt2=-1.857050812e-02 lkt2=-9.991238073e-8 at=1.699105100e+05 lat=-1.189282556e-1 ute=-8.067754816e-01 lute=-2.359536591e-6 ua1=2.393051059e-09 lua1=-7.214822268e-15 pua1=-6.617444900e-36 ub1=-1.688432655e-18 lub1=5.073082956e-24 uc1=-1.199775089e-11 luc1=2.533349999e-16 puc1=-1.033975766e-37 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.165 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.083873259e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.901279921e-9 k1=5.219899191e-01 lk1=1.618360153e-7 k2=-2.203707193e-02 lk2=-7.439951279e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.115866859e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.822597657e-9 nfactor=2.799267766e+00 lnfactor=8.454546788e-7 eta0=0.08 etab=-0.07 u0=2.863473400e-02 lu0=-1.964346373e-9 ua=-4.934718209e-10 lua=-4.578253768e-16 ub=1.172208475e-18 lub=3.122917863e-25 uc=-5.151270940e-12 luc=1.000048738e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.281137600e+04 lvsat=2.671511067e-1 a0=8.439375600e-01 la0=1.296468606e-6 ags=4.376838709e-01 lags=-3.345674742e-7 a1=0.0 a2=0.42385546 b0=2.529228706e-08 lb0=-8.445864377e-14 wb0=6.617444900e-30 b1=3.433965944e-09 lb1=9.339681263e-15 keta=-1.282833575e-02 lketa=6.077299522e-08 wketa=3.469446952e-24 pketa=-2.081668171e-29 dwg=0.0 dwb=0.0 pclm=-7.522176873e-01 lpclm=5.038391298e-6 pdiblc1=0.39 pdiblc2=-6.386343217e-04 lpdiblc2=2.777244603e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.056879617e-01 lkt1=-3.225456744e-8 kt2=-5.679713785e-02 lkt2=5.208189791e-8 at=140000.0 ute=-1.613029847e+00 lute=8.462404173e-7 ua1=-3.252460382e-10 lua1=3.593496680e-15 ub1=6.117920260e-20 lub1=-1.883611737e-24 uc1=5.812970886e-11 luc1=-2.550131747e-17 wuc1=-5.169878828e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.166 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.938526700e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.362373658e-8 k1=6.217111102e-01 lk1=-3.522662043e-8 k2=-6.408281072e-02 lk2=8.688585288e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.797451904e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.107689539e-8 nfactor=3.161729441e+00 lnfactor=1.291811149e-7 eta0=1.556200357e-01 leta0=-1.494354750e-7 etab=-1.380244775e-01 letab=1.344256189e-7 u0=3.175960347e-02 lu0=-8.139513419e-9 ua=-2.373880505e-10 lua=-9.638817346e-16 ub=9.359201014e-19 lub=7.792297471e-25 uc=4.829946030e-11 luc=-5.621040407e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.206681920e+05 lvsat=5.401136973e-2 a0=1.5 ags=3.329123510e-01 lags=-1.275247019e-7 a1=0.0 a2=0.42385546 b0=1.913797268e-07 lb0=-4.126700125e-13 wb0=5.293955920e-29 pb0=7.940933881e-35 b1=1.129183952e-08 lb1=-6.188545585e-15 keta=1.805323083e-02 lketa=-2.531802246e-10 dwg=0.0 dwb=0.0 pclm=2.541215632e+00 lpclm=-1.469880848e-6 pdiblc1=1.953531031e-01 lpdiblc1=3.846487403e-7 pdiblc2=2.081142567e-02 lpdiblc2=-1.461578972e-8 pdiblcb=-0.025 drout=4.680248349e-01 ldrout=1.817554350e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.474223732e-01 lkt1=5.021830556e-8 kt2=-3.432961298e-02 lkt2=7.683013180e-9 at=1.497613600e+05 lat=-1.928977490e-2 ute=-1.639359155e+00 lute=8.982707095e-7 ua1=8.087803889e-10 lua1=1.352506233e-15 ub1=-4.323953449e-19 lub1=-9.082413048e-25 uc1=4.294397687e-11 luc1=4.507754196e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.167 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.158135818e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.218690006e-8 k1=5.952653582e-01 lk1=-9.411969933e-9 k2=-6.385444640e-02 lk2=8.465670656e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.169351653e-01 ldsub=4.203713551e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.066672992e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.259155975e-8 nfactor=3.098600874e+00 lnfactor=1.908031822e-7 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=-1.630640067e-22 peta0=5.898059818e-29 etab=-0.0003125 u0=2.334080442e-02 lu0=7.837940144e-11 ua=-1.285657146e-09 lua=5.937146704e-17 ub=1.885211294e-18 lub=-1.474075602e-25 uc=7.885796353e-11 luc=-3.545029551e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.730898568e+05 lvsat=2.840695574e-3 a0=1.5 ags=3.762869949e-01 lags=-1.698642534e-7 a1=0.0 a2=0.42385546 b0=-4.517147431e-07 lb0=2.150776509e-13 b1=9.667650944e-09 lb1=-4.603116650e-15 keta=3.640521038e-02 lketa=-1.816720814e-8 dwg=0.0 dwb=0.0 pclm=1.429863183e+00 lpclm=-3.850497131e-7 pdiblc1=6.748458678e-01 lpdiblc1=-8.340140914e-8 pdiblc2=1.013619654e-02 lpdiblc2=-4.195314257e-9 pdiblcb=-0.025 drout=3.249506503e-01 ldrout=3.214152972e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.127950400e-07 lalpha0=5.298417792e-13 walpha0=1.588186776e-28 palpha0=-1.588186776e-34 alpha1=0.85 beta0=1.220304672e+01 lbeta0=1.617411747e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.866014421e-01 lkt1=-9.151194823e-9 kt2=-4.153609621e-03 lkt2=-2.177287003e-8 at=2.537953600e+05 lat=-1.208411075e-1 ute=9.716893932e-03 lute=-7.114517882e-7 ua1=3.923378182e-09 lua1=-1.687764798e-15 ub1=-2.711103396e-18 lub1=1.316087658e-24 uc1=-8.391965094e-12 luc1=5.461861525e-17 puc1=-2.584939414e-38 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.168 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='-1.894392775e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.479831754e-07 wvth0=2.833711895e-07 pvth0=-1.349232247e-13 k1=2.755733053e-01 lk1=1.428049254e-07 wk1=-5.312266183e-16 pk1=2.529363385e-22 k2=1.507825200e-02 lk2=-2.911702863e-08 wk2=9.317799864e-09 pk2=-4.436539956e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.890254365e+00 ldsub=-7.546903751e-07 wdsub=-6.486327557e-07 pdsub=3.088374058e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413326e-03 lcdscd=-1.441936607e-09 wcdscd=-4.822274524e-18 pcdscd=2.296059176e-24 cit=0.0 voff='-3.953842317e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=1.248769656e-07 wvoff=1.141295068e-07 pvoff=-5.434116687e-14 nfactor=-8.495759660e+00 lnfactor=5.711295629e-06 wnfactor=4.916879871e-06 pnfactor=-2.341103514e-12 eta0=9.253513184e-01 leta0=-2.072863913e-07 weta0=2.727086470e-09 peta0=-1.298464043e-15 etab=3.920295698e-02 letab=-1.881473162e-08 wetab=-2.293703942e-17 petab=1.092114778e-23 u0=-2.507690271e-03 lu0=1.238577827e-08 wu0=8.745738183e-09 pu0=-4.164160796e-15 ua=-1.064517984e-09 lua=-4.592084904e-17 wua=-3.212126641e-17 pua=1.529409130e-23 ub=2.920531487e-18 lub=-6.403607759e-25 wub=-5.788939296e-25 pub=2.756322401e-31 uc=-8.683275570e-11 luc=4.344102078e-17 wuc=4.325528016e-18 puc=-2.059539608e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=2.400705953e+05 lvsat=-2.905124535e-02 wvsat=-2.260982125e-02 pvsat=1.076534985e-8 a0=1.500000005e+00 la0=-2.231342222e-15 wa0=-1.622799672e-15 pa0=7.726734808e-22 ags=-1.093481874e+00 lags=5.299456168e-07 wags=-3.474567301e-16 pags=1.654362758e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=2.261106420e-01 lketa=-1.084927935e-07 wketa=-5.803514877e-08 pketa=2.763262359e-14 dwg=0.0 dwb=0.0 pclm=3.677243673e-01 lpclm=1.206728138e-07 wpclm=2.255874795e-07 ppclm=-1.074103202e-13 pdiblc1=6.287709947e-01 lpdiblc1=-6.146350335e-08 wpdiblc1=2.778195451e-16 ppdiblc1=-1.322800758e-22 pdiblc2=-5.080122972e-03 lpdiblc2=3.049723249e-09 wpdiblc2=-7.448985873e-18 ppdiblc2=3.546732786e-24 pdiblcb=4.582196904e-02 lpdiblcb=-3.372088905e-08 wpdiblcb=-2.205591265e-17 ppdiblcb=1.050159959e-23 drout=1.449262894e+00 ldrout=-2.139102373e-07 wdrout=-1.471450517e-15 pdrout=7.006102365e-22 pscbe1=8.077610965e+08 lpscbe1=-3.695337436e+00 wpscbe1=-1.453666687e-07 ppscbe1=6.921434402e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.436415553e-06 lalpha0=-3.982475555e-13 walpha0=-1.178617961e-13 palpha0=5.611824414e-20 alpha1=0.85 beta0=1.759308914e+01 lbeta0=-9.489814890e-07 wbeta0=-3.142981258e-07 pbeta0=1.496486524e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.556720410e-01 lkt1=-7.149139618e-08 wkt1=-7.857453133e-08 pkt1=3.741216305e-14 kt2=-6.887994138e-02 lkt2=9.045666669e-09 wkt2=-8.817280239e-18 pkt2=4.198211223e-24 at=1.306347085e+05 lat=-6.219988757e-02 wat=-5.893089846e-02 pat=2.805912227e-8 ute=-1.216531881e+00 lute=-1.275906013e-07 wute=-1.571490625e-07 pute=7.482432602e-14 ua1=7.427581515e-10 lua1=-1.733570997e-16 wua1=-1.663665766e-24 pua1=7.921313156e-31 ub1=-5.392589525e-19 lub1=2.819943316e-25 wub1=-2.363318072e-33 pub1=1.125260585e-39 uc1=6.935515480e-11 luc1=1.760041257e-17 wuc1=3.421922117e-26 puc1=-1.629297653e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.169 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='3.367289995e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.563213553e-07 wvth0=-1.012039962e-06 pvth0=1.580158716e-13 k1=9.070734845e-01 lk1=8.554508213e-16 wk1=1.897239699e-15 pk1=-2.962274870e-22 k2=-4.732794818e-02 lk2=-1.500474014e-08 wk2=-3.327785666e-08 pk2=5.195871427e-15 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=-6.066036018e+00 ldsub=1.044513307e-06 wdsub=2.316545556e-06 pdsub=-3.616961569e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=2.051999950e-03 lcdscd=7.765460150e-18 wcdscd=1.722241447e-17 pcdscd=-2.689038228e-24 cit=0.0 voff='9.695608727e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.837862605e-07 wvoff=-4.076053816e-07 pvoff=6.364187386e-14 nfactor=5.177371864e+01 lnfactor=-7.917803115e-06 wnfactor=-1.756028525e-05 pnfactor=2.741792698e-12 eta0=2.812619630e-02 leta0=-4.391511347e-09 weta0=-9.739594534e-09 peta0=1.520701332e-15 etab=-4.399800024e-02 letab=3.693628736e-17 wetab=8.191813894e-17 petab=-1.279036599e-23 u0=1.145427125e-01 lu0=-1.408353160e-08 wu0=-3.123477923e-08 pu0=4.876873489e-15 ua=-1.496323242e-09 lua=5.172586476e-17 wua=1.147188086e-16 pua=-1.791173590e-23 ub=-4.033564733e-18 lub=9.322107271e-25 wub=2.067478320e-24 pub=-3.228077950e-31 uc=1.360709473e-10 luc=-6.965531008e-18 wuc=-1.544831434e-17 puc=2.412038008e-24 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=-4.940360154e+04 lvsat=3.640929163e-02 wvsat=8.074936160e-02 pvsat=-1.260788232e-8 a0=1.499999983e+00 la0=2.613244732e-15 wa0=5.795715907e-15 pa0=-9.049196947e-22 ags=1.249999996e+00 lags=5.595195418e-16 wags=1.240916703e-15 pags=-1.937512373e-22 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-6.669297466e-01 lketa=9.345578777e-08 wketa=2.072683885e-07 pketa=-3.236205710e-14 dwg=0.0 dwb=0.0 pclm=2.507778499e+00 lpclm=-3.632704673e-07 wpclm=-8.056695698e-07 ppclm=1.257940240e-13 pdiblc1=3.569721529e-01 lpdiblc1=-4.473816873e-16 wpdiblc1=-9.922134225e-16 ppdiblc1=1.549202988e-22 pdiblc2=8.406112023e-03 lpdiblc2=1.199532834e-17 wpdiblc2=2.660351106e-17 ppdiblc2=-4.153767608e-24 pdiblcb=-1.032957702e-01 lpdiblcb=3.551725580e-17 wpdiblcb=7.877121178e-17 ppdiblcb=-1.229899516e-23 drout=5.033266448e-01 ldrout=2.369521024e-15 wdrout=5.255178515e-15 pdrout=-8.205225388e-22 pscbe1=7.914198785e+08 lpscbe1=2.340879440e-07 wpscbe1=5.191669464e-07 ppscbe1=-8.106064796e-14 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-1.163984368e-06 lalpha0=1.897964808e-13 walpha0=4.209349860e-13 palpha0=-6.572310497e-20 alpha1=0.85 beta0=1.115844166e+01 lbeta0=5.061239535e-07 wbeta0=1.122493306e-06 pbeta0=-1.752616149e-13 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.031350325e+00 lkt1=1.265309882e-07 wkt1=2.806233262e-07 pkt1=-4.381540366e-14 kt2=-2.887893909e-02 lkt2=1.419867002e-17 wkt2=3.149014383e-17 pkt2=-4.916747565e-24 at=-5.640717012e+05 lat=9.489824110e-02 wat=2.104674945e-01 pat=-3.286155272e-8 ute=-2.899822368e+00 lute=2.530619761e-07 wute=5.612466518e-07 pute=-8.763080722e-14 ua1=-2.384735316e-11 lua1=2.679052638e-24 wua1=5.941664344e-24 pua1=-9.277077044e-31 ub1=7.077531456e-19 lub1=3.805723081e-33 wub1=8.440420337e-33 pub1=-1.317853387e-39 uc1=1.471862504e-10 luc1=-5.510429087e-26 wuc1=-1.222117996e-25 puc1=1.908160917e-32 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.170 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.9e-07 wmax=4.2e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='-1.552765479e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.118764262e-07 wvth0=8.136238717e-07 pvth0=-1.270359768e-13 k1=0.90707349 k2=-6.861111273e-01 lk2=8.473231032e-08 wk2=1.957465773e-07 pk2=-3.056308759e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.327233918e+00 ldsub=-4.221142877e-07 wdsub=-1.017279861e-06 pdsub=1.588340084e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-9.376860080e+00 lnfactor=1.630003644e-06 wnfactor=1.905910194e-06 pnfactor=-2.975811940e-13 eta0=0.0 etab=-0.043998 u0=2.328525708e-01 lu0=-3.255595964e-08 wu0=-8.966650519e-08 pu0=1.400016945e-14 ua=-1.393966080e-09 lua=3.574422705e-17 wua=1.398486939e-16 pua=-2.183541567e-23 ub=6.496925019e-18 lub=-7.119778210e-25 wub=-2.980183497e-24 pub=4.653139304e-31 uc=-1.261952878e-10 luc=3.398366988e-17 wuc=1.186133762e-16 puc=-1.851981810e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.844848871e+05 lvsat=-3.133632143e-02 wvsat=-9.060217712e-02 pvsat=1.414626153e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.038255850e+00 lketa=1.514331602e-07 wketa=4.029564649e-07 pketa=-6.291601060e-14 dwg=0.0 dwb=0.0 pclm=1.737606982e-02 lpclm=2.557100636e-08 wpclm=1.207637141e-07 ppclm=-1.885556327e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.424179121e-07 lalpha0=-1.417994553e-14 walpha0=2.955654554e-21 palpha0=-4.614840902e-28 alpha1=0.85 beta0=1.671249328e+01 lbeta0=-3.610634506e-07 wbeta0=2.044754410e-14 pbeta0=-3.192596409e-21 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.368700706e-01 lkt1=-1.312958075e-08 wkt1=-1.018287676e-15 pkt1=1.589913756e-22 kt2=-0.028878939 at=1.675154536e+03 lat=6.564790030e-03 wat=-3.270385787e-10 pat=5.106249591e-17 ute=-9.418347041e-01 lute=-5.265038572e-08 wute=-2.218109000e-07 pute=3.463266668e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.171 nmos lmin=2.0e-05 lmax=0.0001 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.4888923+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.56800772 k2=-0.036474946 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=3.3453 eta0=0.08 etab=-0.07 u0=0.0243621 ua=-1.0538187e-9 ub=1.5967e-18 uc=4.8537e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.3626 ags=0.34488 a1=0.0 a2=0.42385546 b0=2.3328e-8 b1=3.9114e-9 keta=-0.0045466 dwg=0.0 dwb=0.0 pclm=0.016875 pdiblc1=0.39 pdiblc2=0.00096032746 pdiblcb=-0.025 drout=0.56 pscbe1=225000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.28638 kt2=-0.029517931 at=175000.0 ute=-1.1154 ua1=1.121e-9 ub1=-5.6947e-19 uc1=3.3818362e-11 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.172 nmos lmin=8.0e-06 lmax=2.0e-05 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.750925212e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=2.756662574e-7 k1=5.566754387e-01 lk1=2.263751931e-7 k2=-2.793918103e-02 lk2=-1.705116018e-7 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.017610378e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.301805274e-7 nfactor=3.511203629e+00 lnfactor=-3.314113452e-6 eta0=0.08 etab=-0.07 u0=2.317604858e-02 lu0=2.369272453e-8 ua=-1.142103671e-09 lua=1.763592594e-15 wua=8.271806126e-31 ub=1.637803688e-18 lub=-8.210928520e-25 uc=6.331678001e-11 luc=-2.952428955e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.478652779e+00 la0=-2.318286092e-6 ags=3.214434537e-01 lags=4.681716359e-7 a1=0.0 a2=0.42385546 b0=1.263931308e-08 lb0=2.135186635e-13 b1=4.228185535e-09 lb1=-6.328150926e-15 keta=-1.968579909e-03 lketa=-5.149887994e-8 dwg=0.0 dwb=0.0 pclm=-2.742977677e-02 lpclm=8.850382462e-07 ppclm=1.110223025e-28 pdiblc1=0.39 pdiblc2=-1.549079328e-04 lpdiblc2=2.227809388e-8 pdiblcb=-0.025 drout=0.56 pscbe1=-6.611043278e+07 lpscbe1=5.815261596e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.785102125e-01 lkt1=-1.572079458e-07 wkt1=-2.220446049e-22 kt2=-2.846841042e-02 lkt2=-2.096536584e-8 at=1.882935600e+05 lat=-2.655539625e-1 ute=-1.123907878e+00 lute=1.699545360e-7 ua1=8.767308350e-10 lua1=4.879554061e-15 ub1=-2.484770535e-19 lub1=-6.412198755e-24 uc1=4.316007430e-11 luc1=-1.866113153e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.173 nmos lmin=4.0e-06 lmax=8.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.096875978e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))' lvth0=-2.687778576e-10 k1=6.072888189e-01 lk1=-1.773240112e-7 k2=-5.783410041e-02 lk2=6.793434087e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.259947907e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=6.311118168e-8 nfactor=3.179000049e+00 lnfactor=-6.644125212e-7 eta0=0.08 etab=-0.07 u0=2.416419740e-02 lu0=1.581111515e-8 ua=-1.231511291e-09 lua=2.476719931e-15 ub=1.817275000e-18 lub=-2.252580446e-24 uc=3.256440823e-11 luc=-4.995779590e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=80000.0 a0=1.205892612e+00 la0=-1.427139067e-7 ags=4.065813044e-01 lags=-2.108994399e-7 a1=0.0 a2=0.42385546 b0=7.455615358e-08 lb0=-2.803384769e-13 b1=1.100708765e-09 lb1=1.861702913e-14 keta=-1.924158216e-02 lketa=8.627293517e-8 dwg=0.0 dwb=0.0 pclm=-3.453042139e-01 lpclm=3.420447988e-06 wpclm=1.110223025e-22 ppclm=-4.440892099e-28 pdiblc1=0.39 pdiblc2=-1.047655494e-03 lpdiblc2=2.939876984e-8 pdiblcb=-0.025 drout=0.56 pscbe1=5.267617483e+08 lpscbe1=1.086432449e+3 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.827329503e-01 lkt1=-1.235268148e-7 kt2=-1.857050812e-02 lkt2=-9.991238073e-8 at=1.699105100e+05 lat=-1.189282556e-1 ute=-8.067754816e-01 lute=-2.359536591e-6 ua1=2.393051059e-09 lua1=-7.214822268e-15 wua1=1.654361225e-30 ub1=-1.688432655e-18 lub1=5.073082956e-24 uc1=-1.199775089e-11 luc1=2.533349999e-16 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.174 nmos lmin=2.0e-06 lmax=4.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.083873259e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=4.901279921e-9 k1=5.219899191e-01 lk1=1.618360153e-7 k2=-2.203707193e-02 lk2=-7.439951279e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.56 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.115866859e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=5.822597657e-9 nfactor=2.799267766e+00 lnfactor=8.454546788e-7 eta0=0.08 etab=-0.07 u0=2.863473400e-02 lu0=-1.964346373e-9 ua=-4.934718209e-10 lua=-4.578253768e-16 ub=1.172208475e-18 lub=3.122917863e-25 uc=-5.151270940e-12 luc=1.000048738e-16 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.281137600e+04 lvsat=2.671511067e-1 a0=8.439375600e-01 la0=1.296468606e-6 ags=4.376838709e-01 lags=-3.345674742e-7 a1=0.0 a2=0.42385546 b0=2.529228706e-08 lb0=-8.445864377e-14 wb0=-3.308722450e-30 pb0=1.985233470e-35 b1=3.433965944e-09 lb1=9.339681263e-15 keta=-1.282833575e-02 lketa=6.077299522e-08 wketa=3.469446952e-24 dwg=0.0 dwb=0.0 pclm=-7.522176873e-01 lpclm=5.038391298e-6 pdiblc1=0.39 pdiblc2=-6.386343217e-04 lpdiblc2=2.777244603e-8 pdiblcb=-0.025 drout=0.56 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.056879617e-01 lkt1=-3.225456744e-8 kt2=-5.679713785e-02 lkt2=5.208189791e-8 at=140000.0 ute=-1.613029847e+00 lute=8.462404173e-7 ua1=-3.252460382e-10 lua1=3.593496680e-15 ub1=6.117920260e-20 lub1=-1.883611737e-24 uc1=5.812970886e-11 luc1=-2.550131747e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=3.0e-6 sbref=3.0e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.175 nmos lmin=1.0e-06 lmax=2.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='4.938526700e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=3.362373658e-8 k1=6.217111102e-01 lk1=-3.522662043e-8 k2=-6.408281072e-02 lk2=8.688585288e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=8.528408000e-01 ldsub=-5.786932471e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-9.797451904e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-2.107689539e-8 nfactor=3.161729441e+00 lnfactor=1.291811149e-7 eta0=1.556200358e-01 leta0=-1.494354750e-7 etab=-1.380244775e-01 letab=1.344256189e-7 u0=3.175960347e-02 lu0=-8.139513419e-9 ua=-2.373880505e-10 lua=-9.638817346e-16 ub=9.359201014e-19 lub=7.792297471e-25 uc=4.829946030e-11 luc=-5.621040407e-18 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.206681920e+05 lvsat=5.401136973e-2 a0=1.5 ags=3.329123510e-01 lags=-1.275247019e-7 a1=0.0 a2=0.42385546 b0=1.913797268e-07 lb0=-4.126700125e-13 wb0=2.646977960e-29 pb0=-7.940933881e-35 b1=1.129183952e-08 lb1=-6.188545585e-15 wb1=-6.617444900e-30 keta=1.805323083e-02 lketa=-2.531802246e-10 dwg=0.0 dwb=0.0 pclm=2.541215632e+00 lpclm=-1.469880848e-6 pdiblc1=1.953531031e-01 lpdiblc1=3.846487403e-7 pdiblc2=2.081142567e-02 lpdiblc2=-1.461578972e-8 pdiblcb=-0.025 drout=4.680248349e-01 ldrout=1.817554350e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=3.0e-8 alpha1=0.85 beta0=13.86 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.474223732e-01 lkt1=5.021830556e-8 kt2=-3.432961298e-02 lkt2=7.683013180e-9 at=1.497613600e+05 lat=-1.928977490e-2 ute=-1.639359155e+00 lute=8.982707095e-7 ua1=8.087803889e-10 lua1=1.352506233e-15 ub1=-4.323953449e-19 lub1=-9.082413048e-25 uc1=4.294397687e-11 luc1=4.507754196e-18 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=2.75e-6 sbref=2.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.176 nmos lmin=5.0e-07 lmax=1.0e-06 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='5.158135818e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.218690006e-8 k1=5.952653582e-01 lk1=-9.411969933e-9 k2=-6.385444640e-02 lk2=8.465670656e-9 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=2.169351653e-01 ldsub=4.203713551e-8 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.0054 cit=0.0 voff='-1.066672992e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-1.259155975e-8 nfactor=3.098600874e+00 lnfactor=1.908031822e-7 eta0=-4.616715915e-01 leta0=4.531251049e-07 weta0=9.367506770e-23 peta0=-9.887923813e-29 etab=-0.0003125 u0=2.334080442e-02 lu0=7.837940144e-11 ua=-1.285657146e-09 lua=5.937146704e-17 ub=1.885211294e-18 lub=-1.474075602e-25 uc=7.885796353e-11 luc=-3.545029551e-17 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.730898568e+05 lvsat=2.840695574e-3 a0=1.5 ags=3.762869949e-01 lags=-1.698642534e-7 a1=0.0 a2=0.42385546 b0=-4.517147431e-07 lb0=2.150776509e-13 b1=9.667650944e-09 lb1=-4.603116650e-15 keta=3.640521038e-02 lketa=-1.816720814e-08 pketa=-6.938893904e-30 dwg=0.0 dwb=0.0 pclm=1.429863183e+00 lpclm=-3.850497131e-7 pdiblc1=6.748458678e-01 lpdiblc1=-8.340140914e-8 pdiblc2=1.013619654e-02 lpdiblc2=-4.195314257e-09 wpdiblc2=6.938893904e-24 pdiblcb=-0.025 drout=3.249506503e-01 ldrout=3.214152972e-7 pscbe1=800000000.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=-5.127950400e-07 lalpha0=5.298417792e-13 walpha0=7.940933881e-29 alpha1=0.85 beta0=1.220304672e+01 lbeta0=1.617411747e-6 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-2.866014421e-01 lkt1=-9.151194823e-9 kt2=-4.153609621e-03 lkt2=-2.177287003e-8 at=2.537953600e+05 lat=-1.208411075e-1 ute=9.716893932e-03 lute=-7.114517882e-7 ua1=3.923378182e-09 lua1=-1.687764798e-15 ub1=-2.711103396e-18 lub1=1.316087658e-24 uc1=-8.391965094e-12 luc1=5.461861525e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.75e-6 sbref=1.74e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.177 nmos lmin=2.5e-07 lmax=5.0e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='6.288856412e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=-4.165077801e-8 k1=2.755733038e-01 lk1=1.428049261e-7 k2=4.198637850e-02 lk2=-4.192895635e-8 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=1.711988033e-02 ldsub=1.371763860e-7 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=8.428413312e-03 lcdscd=-1.441936601e-9 cit=0.0 voff='-6.579878733e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' lvoff=-3.205052951e-8 nfactor=5.703303159e+00 lnfactor=-1.049389345e-6 eta0=9.332265600e-01 leta0=-2.110361214e-7 etab=3.920295691e-02 letab=-1.881473159e-08 wetab=8.673617380e-25 petab=1.192622390e-30 u0=2.274842522e-02 lu0=3.604324679e-10 ua=-1.157278411e-09 lua=-1.754270060e-18 ub=1.248790162e-18 lub=1.556154518e-25 uc=-7.434141045e-11 luc=3.749344162e-17 wuc=-1.292469707e-32 puc=9.693522803e-39 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=1.747775069e+05 lvsat=2.037144600e-3 a0=1.5 ags=-1.093481875e+00 lags=5.299456173e-07 wags=-8.326672685e-23 pags=3.122502257e-29 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=5.851559299e-02 lketa=-2.869475727e-08 pketa=-8.673617380e-31 dwg=0.0 dwb=0.0 pclm=1.019180347e+00 lpclm=-1.895088305e-7 pdiblc1=6.287709955e-01 lpdiblc1=-6.146350373e-8 pdiblc2=-5.080122993e-03 lpdiblc2=3.049723259e-09 wpdiblc2=1.734723476e-24 ppdiblc2=-8.673617380e-31 pdiblcb=4.582196898e-02 lpdiblcb=-3.372088902e-08 ppdiblcb=6.938893904e-30 drout=1.449262890e+00 ldrout=-2.139102352e-7 pscbe1=8.077610961e+08 lpscbe1=-3.695337236e+0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.096051930e-06 lalpha0=-2.361881816e-13 alpha1=0.85 beta0=1.668545280e+01 lbeta0=-5.168231544e-7 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-3.825811247e-01 lkt1=3.654818732e-8 kt2=-6.887994141e-02 lkt2=9.045666681e-9 at=-3.954710419e+04 lat=1.882980000e-2 ute=-1.670350048e+00 lute=8.848856547e-8 ua1=7.427581467e-10 lua1=-1.733570974e-16 ub1=-5.392589593e-19 lub1=2.819943349e-25 wub1=9.629649722e-41 pub1=-3.611118646e-47 uc1=6.935515490e-11 luc1=1.760041252e-17 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.178 nmos lmin=1.8e-07 lmax=2.5e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='0.444701+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' k1=0.90707349 k2=-0.1434284 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=0.62373 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=1.06278 eta0=0.0 etab=-0.043998 u0=0.0243423 ua=-1.165036e-9 ub=1.93694e-18 uc=9.1459e-11 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=183786.0 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-0.068376 dwg=0.0 dwb=0.0 pclm=0.18115 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=5.16e-8 alpha1=0.85 beta0=14.4 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-0.22096074 kt2=-0.028878939 at=43720.487 ute=-1.2790432 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.1e-6 sbref=1.1e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.model sky130_fd_pr__nfet_01v8__model.179 nmos lmin=1.5e-07 lmax=1.8e-07 wmin=3.6e-07 wmax=3.9e-7 level=54.0 version=4.5 binunit=2.0 mobmod=0.0 capmod=2.0 igcmod=0.0 igbmod=0.0 geomod=0.0 diomod=1.0 rdsmod=0.0 rbodymod=1.0 rgatemod=0.0 permod=1.0 acnqsmod=0.0 trnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 tempmod=0.0 toxe='4.148e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))' toxm=4.148e-9 dtox=0.0 epsrox=3.9 xj=1.5e-7 ngate=1.0e+23 ndep=1.7e+17 nsd=1.0e+20 rsh=1.0 rshg=0.1 wint=2.1859e-8 lint=1.1932e-8 vth0='-2.993931675e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))' lvth0=1.161798869e-07 wvth0=3.796036009e-07 pvth0=-5.926978783e-14 k1=0.90707349 k2=-3.222046665e-01 lk2=2.791341115e-08 wk2=6.973232022e-08 pk2=-1.088772555e-14 k3=2.0 k3b=0.54 w0=0.0 dvt0=0.0 dvt1=0.53 dvt2=-0.032 dvt0w=-3.58 dvt1w=1670600.0 dvt2w=0.068 dsub=3.327233912e+00 ldsub=-4.221142868e-07 wdsub=-1.017279859e-06 pdsub=1.588340081e-13 minv=0.0 voffl=5.8197729e-9 lpe0=1.0325e-7 lpeb=-7.082e-8 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 phin=0.0 cdsc=0.0 cdscb=0.0 cdscd=0.002052 cit=0.0 voff='-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))' nfactor=-9.376859947e+00 lnfactor=1.630003623e-06 wnfactor=1.905910148e-06 pnfactor=-2.975811868e-13 eta0=0.0 etab=-0.043998 u0=8.959275208e-02 lu0=-1.018794459e-08 wu0=-4.005820865e-08 pu0=6.254528466e-15 ua=-1.393966070e-09 lua=3.574422544e-17 wua=1.398486904e-16 pua=-2.183541512e-23 ub=6.496924862e-18 lub=-7.119777965e-25 wub=-2.980183442e-24 pub=4.653139219e-31 uc=-1.261952913e-10 luc=3.398367043e-17 wuc=1.186133774e-16 puc=-1.851981829e-23 ud=0.0 up=0.0 lp=1.0 eu=1.67 vtl=0.0 xn=3.0 vsat=3.102888726e+05 lvsat=-1.975165252e-02 wvsat=-6.490943285e-02 pvsat=1.013469921e-8 a0=1.5 ags=1.25 a1=0.0 a2=0.42385546 b0=0.0 b1=0.0 keta=-1.038255847e+00 lketa=1.514331597e-07 wketa=4.029564638e-07 pketa=-6.291601043e-14 dwg=0.0 dwb=0.0 pclm=1.737607849e-02 lpclm=2.557100501e-08 wpclm=1.207637111e-07 ppclm=-1.885556280e-14 pdiblc1=0.35697215 pdiblc2=0.0084061121 pdiblcb=-0.10329577 drout=0.50332666 pscbe1=791419880.0 pscbe2=1.0e-12 pvag=0.0 delta=0.01 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 lambda=0.0 lc=5.0e-9 rdsw=65.968 rsw=0.0 rdw=0.0 rdswmin=0.0 rdwmin=0.0 rswmin=0.0 prwb=0.0 prwg=0.021507 wr=1.0 alpha0=1.424179200e-07 lalpha0=-1.417994676e-14 walpha0=2.191742220e-22 palpha0=-3.422097810e-29 alpha1=0.85 beta0=1.671249334e+01 lbeta0=-3.610634598e-07 wbeta0=3.836930773e-17 pbeta0=-5.989875262e-24 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 toxref=4.148e-9 dlcig=0.0 aigbacc=1.0 bigbacc=0.0 cigbacc=0.0 nigbacc=0.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=0.0 aigc=0.43 bigc=0.054 cigc=0.075 aigsd=0.43 bigsd=0.054 cigsd=0.075 nigc=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 vfbsdoff=0.0 dlc=9.87908e-9 dwc=0.0 xpart=0.0 cgso=2.449068e-10 cgdo=2.449068e-10 cgbo=1.0e-13 cgdl=0.0 cgsl=0.0 clc=1.0e-7 cle=0.6 cf=1.4067e-12 ckappas=0.6 vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.4037 voffcv=-0.17287 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 ef=0.84 noia=2.5e+42 noib=0.0 noic=0.0 em=41000000.0 ntnoi=1.0 lintnoi=-1.0e-7 af=1.0 kf=0.0 tnoia=15000000.0 tnoib=9900000.0 rnoia=0.94 rnoib=0.26 xl=0.0 xw=0.0 dmcg=0.0 dmdg=0.0 dmcgt=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 jss=0.00275 jsws=6.0e-10 ijthsfwd=0.1 ijthsrev=0.1 bvs=11.7 xjbvs=1.0 pbs=0.729 cjs=0.001339749237 mjs=0.44 pbsws=0.2 cjsws=3.67354204e-11 mjsws=0.0009 pbswgs=0.95578 cjswgs=2.38232788e-10 mjswgs=0.8 tnom=30.0 kt1=-1.368700733e-01 lkt1=-1.312958033e-08 wkt1=-8.156852971e-17 pkt1=1.273581240e-23 kt2=-0.028878939 at=1.675153666e+03 lat=6.564790165e-03 wat=-2.587959170e-11 pat=4.040746717e-18 ute=-9.418347116e-01 lute=-5.265038454e-08 wute=-2.218108973e-07 pute=3.463266627e-14 ua1=-2.3847336e-11 ub1=7.0775317e-19 uc1=1.4718625e-10 kt1l=0.0 prt=0.0 tvoff=0.0 njs=1.2928 tpb=0.0012287 tcj=0.000792 tpbsw=0.0 tcjsw=1.0e-5 tpbswg=0.0 tcjswg=0.0 xtis=2.0 tvfbsdoff=0.0 ll=0.0 wl=0.0 lln=1.0 wln=1.0 lw=0.0 ww=0.0 lwn=1.0 wwn=1.0 lwl=0.0 wwl=0.0 llc=0.0 wlc=0.0 lwc=0.0 wwc=0.0 lwlc=0.0 wwlc=0.0 saref=1.04e-6 sbref=1.04e-6 kvth0=9.8e-9 lkvth0=0.0 wkvth0=2.0e-7 pkvth0=0.0 llodvth=0.0 wlodvth=1.0 wlod=0.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0=-2.7e-8 lku0=0.0 wku0=0.0 pku0=0.0 tku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat=0.2 steta0=0.0
.ends sky130_fd_pr__nfet_01v8