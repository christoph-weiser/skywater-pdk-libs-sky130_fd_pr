* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_bs_flash__special_sonosfet_star__tox_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__ajunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__pjunction_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__overlap_mult=1.0
.param sky130_fd_bs_flash__special_sonosfet_star__lint_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__wint_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__dlc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__dwc_diff=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__k2_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__vth0_diff_0=9.1203e-1
.param sky130_fd_bs_flash__special_sonosfet_star__vsat_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__u0_diff_0=-6.9221e-3
.param sky130_fd_bs_flash__special_sonosfet_star__kt1_diff_0=-4.4275e-1
.param sky130_fd_bs_flash__special_sonosfet_star__nfactor_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__rdsw_diff_0=0.0
.param sky130_fd_bs_flash__special_sonosfet_star__voff_diff_0=0.0