* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__rf_aura_drc_flag_check b_p nwell vgnd
xsky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_1 sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_1/drain sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_1/source sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_1/gate subs sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_0 sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_0/drain sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_0/gate sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_0/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_1 sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_1/drain sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_1/gate sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_1/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_2 sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_2/drain sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_2/gate sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_2/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15
xsky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_0 sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_0/drain sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_0/gate sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_0/source b_p subs sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15
xsky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_1 sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_1/drain sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_2/gate sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_1/source b_p subs sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15
xsky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_3 sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_3/drain sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_3/gate sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_3/source b_p subs sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_0 sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_0/drain sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_0/source sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_1/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15
xsky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_2 sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_2/drain sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_2/gate sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_2/source b_p subs sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_0 sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_0/drain sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_0/gate sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_0/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_1 sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_1/drain sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_1/source sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_1/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_1 sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_1/drain sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_4/gate sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_1/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_2 sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_2/drain sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_3/source sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_2/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_3 sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_3/drain sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_3/source sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15_3/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w0p84l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_2 sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_2/drain sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_2/gate sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_2/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_3 sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_3/drain sky130_fd_pr__rf_nfet_01v8_lvt_af08w3p00l0p15_2/gate sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_3/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_1 sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_1/drain sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_1/source sky130_fd_pr__rf_pfet_01v8_af04w1p68l0p15_3/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_0 sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_0/drain sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_2/source sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_0/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_4 sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_4/drain sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_4/gate sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_4/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
xsky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_2 sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_2/drain sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_2/source sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15_2/gate b_p subs sky130_fd_pr__rf_pfet_01v8_af02w5p00l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_5 sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_5/drain sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_5/gate sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15_5/source subs sky130_fd_pr__rf_nfet_01v8_lvt_af02w0p42l0p15
xsky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_0 sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_0/drain sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_0/source sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15_1/gate subs sky130_fd_pr__rf_nfet_01v8_lvt_af04w0p84l0p15
.ends