* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre=0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre=0.0
.subckt sky130_fd_pr__pfet_01v8_lvt d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param sa=0
.param sb=0
.param sd=0
.param mult=1
.param nf=1.0
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs' sa='sa' sb='sb' sd='sd' nf='nf'
.model sky130_fd_pr__pfet_01v8_lvt__model.0 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-0.29976+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' k1=0.64774 k2=0.002336 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.0054e-9 ub=3.0419e-18 uc=4.9353e-11 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=0.00225131 a0=1.74812 keta=-0.01258 a1=0.0 a2=0.46703705 ags=0.279274 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.154373+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5411305+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=0.0018466 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=0.01363 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.97183 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.1 pmos lmin=8e-06 lmax=2.0e-05 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-0.29976+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' k1=0.64774 k2=0.002336 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.0054e-9 ub=3.0419e-18 uc=4.9353e-11 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=0.00225131 a0=1.74812 keta=-0.01258 a1=0.0 a2=0.46703705 ags=0.279274 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-0.154373+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' nfactor='2.5411305+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=0.0018466 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=0.01363 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-0.97183 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.2 pmos lmin=4e-06 lmax=8e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.029772969e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.560887880e-8 k1=0.64774 k2=-6.558837500e-05 lk2=1.911604307e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.063707319e-09 lua=4.641116804e-16 ub=3.130202425e-18 lub=-7.028652274e-25 uc=3.789249356e-11 luc=9.122276612e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.171669528e-03 lu0=6.339182460e-10 a0=1.837184677e+00 la0=-7.089325618e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.645664986e-01 lags=1.170680346e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.399268421e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.149878056e-7 nfactor='2.472821348e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=5.437237749e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=9.025288750e-05 lpdiblc2=1.398008393e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.927296312e-03 ldelta=6.131159568e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.077060356e+00 lkt1=8.376073282e-7 kt2=-0.055045 at=2.990532506e+05 lat=-1.070845117e-1 ute=-3.115370919e-01 lute=7.070414446e-7 ua1=6.683900700e-10 lua1=1.096847978e-16 ub1=-1.751307275e-19 lub1=2.108595682e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.3 pmos lmin=2e-06 lmax=4e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.610914382e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.402486499e-7 k1=0.64774 k2=-1.116390838e-02 lk2=6.306261569e-08 pk2=-2.524354897e-29 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.561076335e+05 lvsat=-1.280885418e-1 ua=-3.110237112e-09 lua=6.483580312e-16 ub=3.171996025e-18 lub=-8.683574350e-25 uc=6.135820537e-11 luc=-1.695586234e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.033652629e-03 lu0=1.180430663e-9 a0=2.205121124e+00 la0=-2.165868910e-06 wa0=-3.388131789e-21 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.359579442e-01 lags=-1.656242425e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.461535301e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-9.033167759e-8 nfactor='2.607217892e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.154705865e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=3.221488000e-04 lpdiblc2=1.306183409e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.970993700e-02 ldelta=6.735784214e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-9.186784200e-01 lkt1=2.104544561e-7 kt2=-0.055045 at=3.761903100e+05 lat=-4.125279825e-1 ute=-0.13298 ua1=6.9609e-10 ub1=-1.565136819e-19 lub1=1.371407218e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.4 pmos lmin=1.5e-06 lmax=2e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.421589725e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.862345036e-8 k1=0.64774 k2=1.089182255e-01 lk2=-1.722683462e-7 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=90748.0 ua=-2.247467100e-09 lua=-1.042455501e-15 ub=1.852758050e-18 lub=1.717019187e-24 uc=2.825296150e-11 luc=6.318241545e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.934917605e-03 lu0=-5.858233739e-10 a0=1.029745622e+00 la0=1.375732301e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.831765798e-01 lags=1.337890365e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.410403115e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=9.562269231e-8 nfactor='2.576385609e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.197062428e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-3.040698600e-03 lpdiblc2=1.965217428e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.711239350e-02 ldelta=1.182632009e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.096038150e-01 lkt1=-1.992795011e-7 kt2=-0.055045 at=2.048988850e+05 lat=-7.683961238e-2 ute=-0.13298 ua1=7.976886000e-10 lua1=-1.991078563e-16 ub1=-3.072346025e-19 lub1=4.325160460e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.5 pmos lmin=1e-06 lmax=1.5e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.100351645e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.826927837e-8 k1=0.64774 k2=-4.271020350e-02 lk2=4.907125306e-08 pk2=2.524354897e-29 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=9.005122150e+04 lvsat=1.017122415e-3 ua=-3.146447850e-09 lua=2.698316490e-16 ub=3.137067850e-18 lub=-1.577520440e-25 uc=6.944758400e-11 luc=3.048565256e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.825611620e-03 lu0=1.033486038e-9 a0=9.977252900e-01 la0=1.843149104e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-5.337403630e-02 lags=4.790937983e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.519895130e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.436921087e-8 nfactor='2.688930766e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-9.231716865e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=9.396700000e-04 lpdiblc2=1.384183122e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.075824550e-02 ldelta=2.110178763e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.767300750e-01 lkt1=-1.012919430e-7 kt2=-9.202608700e-02 lkt2=5.398314175e-8 at=2.025317050e+05 lat=-7.338412137e-2 ute=4.956445000e-02 lute=-2.664692609e-7 ua1=6.6129e-10 ub1=-1.051962950e-20 lub1=-6.136358374e-28 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.6 pmos lmin=5e-07 lmax=1e-06 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.335619835e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.689413836e-9 k1=0.64774 k2=2.604029800e-02 lk2=-1.691204076e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=9.418488850e+04 lvsat=-2.950164488e-3 ua=-2.795142150e-09 lua=-6.733399654e-17 ub=2.835418650e-18 lub=1.317557757e-25 uc=7.554065400e-11 luc=-2.799258677e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.910283335e-03 lu0=-7.527640766e-12 a0=1.275936345e+00 la0=-8.269814961e-8 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.687461690e-01 lags=-2.201106870e-8 b0=7.194076050e-08 lb0=-6.904514489e-14 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.401774480e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.570584030e-8 nfactor='2.540277169e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=5.035312155e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-2.007644950e-02 lpdiblc2=3.401205191e-08 ppdiblc2=-1.262177448e-29 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.216615250e-02 ldelta=1.015304889e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.147598650e-01 lkt1=-2.567428521e-7 kt2=-1.717199800e-02 lkt2=-1.785807017e-8 at=1.874319130e+05 lat=-5.889209600e-2 ute=-7.139720000e-02 lute=-1.503763173e-7 ua1=4.451523300e-10 lua1=2.074381288e-16 ub1=5.295630895e-19 lub1=-5.189580254e-25 wub1=4.591774808e-41 pub1=3.503246161e-46 uc1=-2.194613080e-11 luc1=1.150272929e-17 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.7 pmos lmin=3.5e-07 lmax=5e-07 wmin=7e-06 wmax=1.0e-4 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.374182550e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=8.803350699e-8 k1=0.64774 k2=-9.546782000e-02 lk2=3.895131649e-08 wk2=5.293955920e-23 pk2=2.524354897e-29 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-5.564831500e+04 lvsat=6.593565082e-2 ua=-3.060750500e-09 lua=5.477944238e-17 ub=3.039400000e-18 lub=3.797535000e-26 uc=8.249041000e-11 luc=-5.994408998e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.709192650e-03 lu0=-3.748261983e-10 a0=1.294423900e+00 la0=-9.119780303e-8 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.120937500e-01 lags=4.034880938e-9 b0=-2.398025350e-07 lb0=7.427883522e-14 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='5.705240200e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.724508402e-07 pvoff=2.019483917e-28 nfactor='-1.363788750e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.488264328e-06 pnfactor=3.231174268e-27 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-7.416210500e-02 lpdiblc2=5.887793202e-8 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.684411500e-02 ldelta=8.002355629e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.456703850e+00 lkt1=1.303408950e-7 kt2=-0.056015 at=1.297958650e+05 lat=-3.239392293e-2 ute=-0.39848 ua1=8.9635e-10 ub1=-5.9922e-19 uc1=3.0734e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.8 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.119795432e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=8.614042311e-8 k1=0.64774 k2=2.404998300e-04 wk2=1.477201471e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.123303443e-09 wua=8.311482974e-16 ub=3.234534534e-18 wub=-1.357957497e-24 uc=5.089054169e-11 wuc=-1.083874332e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.267518568e-03 wu0=-1.142606439e-10 a0=1.722847763e+00 wa0=1.781540569e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.947087473e-01 wags=-1.088056770e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-8.729308566e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-4.728730140e-7 nfactor='2.392497683e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=1.047771884e-6 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.357346608e-03 wpdiblc2=-3.600456115e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.354475070e-03 wdelta=7.243626489e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.560220569e-01 wkt1=-8.163762827e-7 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.9 pmos lmin=8e-06 lmax=2.0e-05 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.119795432e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=8.614042311e-8 k1=0.64774 k2=2.404998300e-04 wk2=1.477201471e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.123303443e-09 wua=8.311482974e-16 ub=3.234534534e-18 wub=-1.357957497e-24 uc=5.089054169e-11 wuc=-1.083874332e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.267518568e-03 wu0=-1.142606439e-10 a0=1.722847763e+00 wa0=1.781540569e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.947087473e-01 wags=-1.088056770e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-8.729308566e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-4.728730140e-7 nfactor='2.392497683e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=1.047771884e-6 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.357346608e-03 wpdiblc2=-3.600456115e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.354475070e-03 wdelta=7.243626489e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.560220569e-01 wkt1=-8.163762827e-7 kt2=-0.055045 at=285600.0 ute=-0.22271 ua1=6.8217e-10 ub1=-1.4864e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.10 pmos lmin=4e-06 lmax=8e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.784072292e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.672272263e-07 wvth0=-1.732041861e-07 pvth0=2.064318253e-12 k1=0.64774 k2=1.829063603e-02 lk2=-1.436745716e-07 wk2=-1.294003316e-07 pk2=1.147575833e-12 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.328819191e-09 lua=1.635853976e-15 wua=1.868879105e-15 pua=-8.260077794e-21 ub=3.545774003e-18 lub=-2.477388364e-24 wub=-2.929529449e-24 pub=1.250931985e-29 uc=1.049570611e-11 luc=3.215327925e-16 wuc=1.931308587e-16 puc=-1.623547039e-21 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.996607109e-03 lu0=2.156387480e-09 wu0=1.234084665e-09 pu0=-1.073249157e-14 a0=2.038498454e+00 la0=-2.512500584e-06 wa0=-1.419140935e-06 pa0=1.271406881e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.280214353e-01 lags=-2.651606682e-07 wags=-4.473191043e-07 pags=2.694482253e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='7.259707909e-04+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.006096846e-07 wvoff=-9.915176576e-07 pvoff=4.128281702e-12 nfactor='2.087826528e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.425106228e-06 wnfactor=2.713981715e-06 pnfactor=-1.326261370e-11 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.080502740e-04 lpdiblc2=1.962394283e-08 wpdiblc2=1.397917910e-09 ppdiblc2=-3.978580764e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-1.202606045e-02 ldelta=1.224252176e-07 wdelta=1.265603573e-07 pdelta=-4.308142442e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.950743407e-01 lkt1=-4.851285840e-07 wkt1=-1.987831654e-06 pkt1=9.324491893e-12 kt2=-0.055045 at=2.990532506e+05 lat=-1.070845117e-1 ute=-3.115370919e-01 lute=7.070414446e-7 ua1=6.683900700e-10 lua1=1.096847978e-16 ub1=-1.751307275e-19 lub1=2.108595682e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.11 pmos lmin=2e-06 lmax=4e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-1.307811179e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-8.517897205e-07 wvth0=-9.186093119e-07 pvth0=5.015936200e-12 k1=0.64774 k2=-7.616810419e-02 lk2=2.303584250e-07 wk2=4.582404480e-07 pk2=-1.179334743e-12 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=2.377756714e+05 lvsat=-4.514735550e-01 wvsat=-5.757105034e-01 pvsat=2.279669666e-6 ua=-3.639276963e-09 lua=2.865189138e-15 wua=3.729412466e-15 pua=-1.562732477e-20 ub=3.986487150e-18 lub=-4.222502247e-24 wub=-5.741672105e-24 pub=2.364470173e-29 uc=1.112943566e-10 luc=-7.760466378e-17 wuc=-3.520198046e-16 puc=5.351132994e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.257701511e-03 lu0=5.082268923e-09 wu0=5.469988258e-09 pu0=-2.750561083e-14 a0=3.343004890e+00 la0=-7.678019947e-06 wa0=-8.021395544e-06 pa0=3.885734650e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.403955315e-01 lags=-7.101339954e-07 wags=-7.362221184e-07 pags=3.838465963e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='4.092964808e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-8.598061957e-07 wvoff=-1.318823782e-06 pvoff=5.424332129e-12 nfactor='2.129443588e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.260313072e-06 wnfactor=3.368021222e-06 pnfactor=-1.585244664e-11 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.444947878e-03 lpdiblc2=9.514708398e-09 wpdiblc2=-1.496445557e-08 ppdiblc2=2.500510075e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.338684151e-02 ldelta=-5.739852094e-08 wdelta=-9.641394332e-08 pdelta=4.521082425e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.084165544e+00 lkt1=6.596003079e-07 wkt1=1.166584600e-06 pkt1=-3.166207869e-12 kt2=-0.055045 at=5.786534212e+05 lat=-1.214231287e+00 wat=-1.427243051e+00 pat=5.651525671e-6 ute=-0.13298 ua1=6.9609e-10 ub1=-2.439533039e-19 lub1=4.833797650e-25 wub1=6.163966964e-25 pub1=-2.440776819e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.12 pmos lmin=1.5e-06 lmax=2e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-9.432847866e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=7.405143442e-07 wvth0=4.237575111e-06 pvth0=-5.088896223e-12 k1=0.64774 k2=2.901341730e-01 lk2=-4.875024628e-07 wk2=-1.277463338e-06 pk2=2.222210751e-12 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-3.845648890e+05 lvsat=7.681583582e-01 wvsat=3.350669729e+00 pvsat=-5.415053994e-6 ua=-5.072658005e-10 lua=-3.272769738e-15 wua=-1.226737156e-14 pua=1.572237272e-20 ub=-7.882126803e-19 lub=5.134715744e-24 wub=1.861725378e-23 pub=-2.409270328e-29 uc=5.379137119e-11 luc=3.508681188e-17 wuc=-1.800304142e-16 puc=1.980570916e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=6.166400069e-03 lu0=-4.537553075e-09 wu0=-2.278000602e-08 pu0=2.785731545e-14 a0=-1.068396601e+00 la0=9.672241253e-07 wa0=1.479063959e-05 pa0=-5.848539361e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=8.662496201e-01 lags=-1.544701546e-06 wags=-4.815253724e-06 pags=1.183234815e-11 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-8.300202179e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=8.470378042e-07 wvoff=4.151953774e-06 pvoff=-5.297024187e-12 nfactor='4.076959946e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.556332109e-06 wnfactor=-1.057814573e-05 pnfactor=1.147855403e-11 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-6.473021715e-03 lpdiblc2=2.699169931e-08 wpdiblc2=2.419581170e-08 ppdiblc2=-5.173923304e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-6.447425998e-03 ldelta=2.066668481e-08 wdelta=1.660825445e-07 pdelta=-6.231924940e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-4.000875206e-01 lkt1=-6.810215983e-07 wkt1=-2.181903547e-06 pkt1=3.395991777e-12 kt2=-2.051672798e-01 lkt2=2.942021378e-07 wkt2=1.058271699e-06 pkt2=-2.073947962e-12 at=-8.405999133e+05 lat=1.567150435e+00 wat=7.370137138e+00 pat=-1.158914015e-5 ute=-0.13298 ua1=8.435353413e-10 lua1=-2.889560076e-16 wua1=-3.231919265e-16 pua1=6.333753779e-22 ub1=4.252388548e-20 lub1=-7.804390684e-26 wub1=-2.465586786e-24 pub1=3.599140310e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.13 pmos lmin=1e-06 lmax=1.5e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-5.152352930e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.156690960e-07 wvth0=1.446537376e-06 pvth0=-1.014678888e-12 k1=0.64774 k2=-1.834256795e-01 lk2=2.037765319e-07 wk2=9.919593950e-07 pk2=-1.090579083e-12 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=4.190611777e+05 lvsat=-4.049347925e-01 wvsat=-2.319322127e+00 pvsat=2.861716617e-6 ua=-3.206959457e-09 lua=6.681080769e-16 wua=4.265704008e-16 pua=-2.807609054e-21 ub=3.110224872e-18 lub=-5.560284719e-25 wub=1.892268388e-25 pub=2.807609054e-30 uc=1.035560908e-10 luc=-3.755723751e-17 wuc=-2.404444393e-16 puc=2.862464648e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.815580322e-03 lu0=1.813556050e-09 wu0=7.071461327e-11 pu0=-5.499023985e-15 a0=-1.788868640e+00 la0=2.018933184e-06 wa0=1.964380967e-05 pa0=-1.293295439e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-1.533070986e+00 lags=1.957706709e-06 wags=1.043097272e-05 pags=-1.042333090e-11 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.962752918e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=6.790364832e-08 wvoff=1.017127881e-06 pvoff=-7.209620890e-13 nfactor='3.777138492e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.118667742e-06 wnfactor=-7.671209360e-06 pnfactor=7.235153676e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.741299014e-02 lpdiblc2=-7.875906499e-09 wpdiblc2=-1.161269901e-07 ppdiblc2=1.530969768e-13 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.520137611e-03 ldelta=3.197033833e-09 wdelta=3.692550728e-08 pdelta=1.262177356e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.898644681e-01 lkt1=-1.120446992e-07 wkt1=9.258956438e-08 pkt1=7.580045758e-14 kt2=5.809619276e-02 lkt2=-9.009671626e-08 wkt2=-1.058271699e-06 pkt2=1.015676263e-12 at=9.217763381e+05 lat=-1.005478298e+00 wat=-5.070241678e+00 pat=6.570702823e-6 ute=3.300117136e-01 lute=-6.758521539e-07 wute=-1.976984379e-06 pute=2.885902947e-12 ua1=5.192954496e-10 lua1=1.843531742e-16 wua1=1.000976099e-15 pua1=-1.299578898e-21 ub1=-9.458320519e-21 lub1=-2.162881622e-27 wub1=-7.481589408e-27 pub1=1.092125014e-32 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.14 pmos lmin=5e-07 lmax=1e-06 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.369118879e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-5.547679202e-08 wvth0=2.361480968e-08 pvth0=3.509710442e-13 k1=0.64774 k2=6.047475350e-02 lk2=-3.030690864e-08 wk2=-2.427421817e-07 pk2=9.442575484e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=7.831437685e+04 lvsat=-7.790305044e-02 wvsat=1.118775531e-01 pvsat=5.283727243e-7 ua=-1.814808597e-09 lua=-6.680087105e-16 wua=-6.910761385e-15 pua=4.234395127e-21 ub=1.545566720e-18 lub=9.456521889e-25 wub=9.092679615e-24 pub=-5.737479748e-30 uc=3.800181094e-11 luc=2.535848255e-17 wuc=2.646262452e-16 puc=-1.984951247e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.471759640e-03 lu0=-7.357120501e-10 wu0=-1.100746794e-08 pu0=5.133261719e-15 a0=1.151289885e+00 la0=-8.028839602e-07 wa0=8.786825050e-07 pa0=5.076876413e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.998143349e-01 lags=1.026200224e-07 wags=4.859279333e-07 pags=-8.785741641e-13 b0=1.276335481e-06 lb0=-1.224962978e-12 wb0=-8.490257731e-12 pb0=8.148524858e-18 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.296030253e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-9.206005949e-08 wvoff=-7.454331392e-08 pvoff=3.267693400e-13 nfactor='2.498382706e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.086181232e-07 wnfactor=2.953307410e-07 pnfactor=-4.107331861e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-3.820576011e-02 lpdiblc2=4.550418905e-08 wpdiblc2=1.278007260e-07 ppdiblc2=-8.101264862e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=4.231590859e-03 ldelta=4.433716578e-09 wdelta=1.264278630e-07 pdelta=4.031784975e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.530963716e-01 lkt1=-2.433078798e-07 wkt1=2.702492927e-07 pkt1=-9.470846668e-14 kt2=-1.717199800e-02 lkt2=-1.785807017e-8 at=-2.961663665e+05 lat=1.634422130e-01 wat=3.409076744e+00 pat=-1.567323033e-6 ute=-3.518444636e-01 lute=-2.144068786e-08 wute=1.976984379e-06 pute=-9.089185683e-13 ua1=5.413001391e-10 lua1=1.632341736e-16 wua1=-6.777841728e-16 pua1=3.116112735e-22 ub1=5.285017805e-19 lub1=-5.184700886e-25 wub1=7.481589408e-27 pub1=-3.439660730e-33 uc1=-2.194613080e-11 luc1=1.150272929e-17 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.15 pmos lmin=3.5e-07 lmax=5e-07 wmin=5.0e-06 wmax=7.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-8.815305629e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.949116438e-07 wvth0=2.425784615e-06 pvth0=-7.534265240e-13 k1=0.64774 k2=-1.109182205e-01 lk2=4.849101115e-08 wk2=1.089160222e-07 pk2=-6.724910441e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-8.773932710e+05 lvsat=3.614835407e-01 wvsat=5.792807249e+00 pvsat=-2.083434704e-6 ua=-4.060526255e-09 lua=3.644599824e-16 wua=7.047817205e-15 pua=-2.183061379e-21 ub=4.511979923e-18 lub=-4.181562813e-25 wub=-1.038080197e-23 pub=3.215453409e-30 uc=1.551521309e-10 luc=-2.850137704e-17 wuc=-5.122213897e-16 puc=1.586605755e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.596554919e-03 lu0=-7.930866800e-10 wu0=-6.255369806e-09 pu0=2.948484603e-15 a0=-3.888856237e+00 la0=1.514323219e-06 wa0=3.653900463e-05 pa0=-1.131795668e-11 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.054057549e+00 lags=-1.981682952e-07 wags=-4.525458319e-06 pags=1.425410665e-12 b0=-4.254451602e-06 lb0=1.317816384e-12 wb0=2.830085910e-11 pb0=-8.766191108e-18 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='2.939064976e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.867685626e-07 wvoff=1.949987009e-06 pvoff=-6.040084762e-13 nfactor='-1.337786068e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.407721022e-06 wnfactor=-1.833032520e-06 pnfactor=5.677818230e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.364520468e-01 lpdiblc2=9.067291935e-08 wpdiblc2=4.391065910e-07 ppdiblc2=-2.241355201e-13 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.407641743e-03 ldelta=5.272277184e-09 wdelta=1.722624257e-07 pdelta=1.924540953e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.581766330e+00 lkt1=1.836481335e-07 wkt1=8.816151949e-07 pkt1=-3.757839402e-13 kt2=-0.056015 at=1.297958650e+05 lat=-3.239392293e-2 ute=-0.39848 ua1=8.9635e-10 ub1=-5.9922e-19 uc1=3.0734e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.16 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.931665961e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=-8.853633893e-9 k1=0.64774 k2=1.017046721e-02 wk2=-3.536834270e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.111169900e-09 wua=7.698812081e-16 ub=3.072328930e-18 wub=-5.389168457e-25 uc=3.016401799e-11 wuc=9.381772402e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.905370027e-03 wu0=1.714371474e-9 a0=1.760051121e+00 wa0=-9.700503222e-9 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.899405748e-01 wags=-8.472927636e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.785927869e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-1.186448532e-8 nfactor='2.581383901e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=9.401019432e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=7.244490933e-04 wpdiblc2=4.644693329e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.317621807e-02 wdelta=2.284237544e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.151583819e+00 wkt1=6.760326889e-7 kt2=-0.055045 at=2.899606391e+05 wat=-2.201860255e-2 ute=-1.174447810e-01 wute=-5.315259861e-7 ua1=6.8217e-10 ub1=-1.463681985e-19 wub1=-1.147123000e-26 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.17 pmos lmin=8e-06 lmax=2.0e-05 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.931665962e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=-8.853633893e-9 k1=0.64774 k2=1.017046721e-02 wk2=-3.536834270e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.111169900e-09 wua=7.698812081e-16 ub=3.072328930e-18 wub=-5.389168457e-25 uc=3.016401799e-11 wuc=9.381772402e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.905370027e-03 wu0=1.714371474e-9 a0=1.760051121e+00 wa0=-9.700503222e-9 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.899405748e-01 wags=-8.472927636e-8 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.785927869e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-1.186448532e-8 nfactor='2.581383901e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=9.401019432e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=7.244490933e-04 wpdiblc2=4.644693329e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.317621807e-02 wdelta=2.284237544e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.151583819e+00 wkt1=6.760326889e-7 kt2=-0.055045 at=2.899606391e+05 wat=-2.201860255e-2 ute=-1.174447810e-01 wute=-5.315259861e-7 ua1=6.8217e-10 ub1=-1.463681985e-19 wub1=-1.147123000e-26 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.18 pmos lmin=4e-06 lmax=8e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.963452000e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.530089208e-08 wvth0=-8.262823205e-08 pvth0=5.872273577e-13 k1=0.64774 k2=-9.174101374e-04 lk2=8.825673168e-08 wk2=-3.241126170e-08 pk2=-2.353762549e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.156450601e-09 lua=3.604230637e-16 wua=9.985214917e-16 pua=-1.819919497e-21 ub=3.072328930e-18 wub=-5.389168457e-25 uc=3.016401799e-11 wuc=9.381772402e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.723853280e-03 lu0=1.444827926e-09 wu0=2.611327307e-09 pu0=-7.139544186e-15 a0=1.847722787e+00 la0=-6.978445481e-07 wa0=-4.558386671e-07 pa0=3.551148250e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.391096336e-01 lags=4.046015844e-07 wags=1.631969404e-09 pags=-6.874139260e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.937541549e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=1.206806989e-07 wvoff=-9.510100109e-09 pvoff=-1.874031770e-14 nfactor='2.562835735e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.476387600e-07 wnfactor=3.154711730e-07 pnfactor=-1.762774025e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.513579764e-03 lpdiblc2=1.781415019e-08 wpdiblc2=8.494995703e-09 ppdiblc2=-3.064744433e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.180500002e-02 ldelta=1.091455284e-08 wdelta=6.227848174e-09 pdelta=1.322474834e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.455881131e+00 lkt1=2.422130526e-06 wkt1=1.348844830e-06 pkt1=-5.355416440e-12 kt2=-0.055045 at=3.077306500e+05 lat=-1.414448437e-01 wat=-4.381564292e-02 pat=1.734989920e-7 ute=-1.020658852e-01 lute=-1.224121660e-07 wute=-1.057703492e-06 pute=4.188241402e-12 ua1=6.683900700e-10 lua1=1.096847978e-16 ub1=-1.706099845e-19 lub1=1.929585561e-25 wub1=-2.282703075e-26 pub1=9.038933501e-32 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.19 pmos lmin=2e-06 lmax=4e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.635397667e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=2.913745773e-07 wvth0=2.566817438e-07 pvth0=-7.563553191e-13 k1=0.64774 k2=2.008035702e-02 lk2=5.110823202e-09 wk2=-2.775633954e-08 pk2=-4.196995353e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.918974676e-09 lua=-5.799222339e-16 wua=9.231953519e-17 pua=1.768413700e-21 ub=2.778925643e-18 lub=1.161803665e-24 wub=3.557865500e-25 pub=-3.542801771e-30 uc=-2.490208249e-12 luc=1.293025723e-16 wuc=2.225237496e-16 puc=-5.096436848e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.281704706e-03 lu0=-7.641242571e-10 wu0=2.993885749e-10 pu0=2.015155206e-15 a0=1.362747454e+00 la0=1.222536528e-06 wa0=1.977712395e-06 pa0=-6.085105568e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.992914103e-01 lags=1.662967941e-07 wags=-2.373125142e-08 pags=-5.869819123e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.491668848e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=3.401012562e-07 wvoff=1.459890705e-07 pvoff=-6.344781587e-13 nfactor='3.096892361e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.967091965e-06 wnfactor=-1.517012678e-06 pnfactor=5.493403903e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.408670462e-03 lpdiblc2=1.739873559e-08 wpdiblc2=4.493997166e-09 ppdiblc2=-1.480449037e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.266166368e-02 ldelta=7.522378933e-09 wdelta=8.235728198e-09 pdelta=1.242967805e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.502781021e-01 lkt1=2.409393284e-08 wkt1=-1.440618077e-08 pkt1=4.271674985e-14 kt2=-0.055045 at=2.848968128e+05 lat=-5.102855685e-02 wat=5.605098002e-02 pat=-2.219478681e-7 ute=-0.13298 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.20 pmos lmin=1.5e-06 lmax=2e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='7.387640686e-03+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-4.355504092e-07 wvth0=-5.627483414e-07 pvth0=8.495227903e-13 k1=0.64774 k2=4.209401888e-02 lk2=-3.803045063e-08 wk2=-2.500987975e-08 pk2=-4.735232809e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=5.157275256e+05 lvsat=-7.681583582e-01 wvsat=-1.195264989e+00 pvsat=2.342420561e-6 ua=-3.009981238e-09 lua=-4.015721230e-16 wua=3.698347649e-16 pua=1.224553229e-21 ub=2.903708702e-18 lub=9.172600652e-25 wub=-2.472665970e-26 pub=-2.797091008e-30 uc=-3.224380557e-11 luc=1.876121847e-16 wuc=2.543954352e-16 puc=-5.721042207e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=8.850258880e-04 lu0=1.973017056e-09 wu0=3.887754209e-09 pu0=-5.017144344e-15 a0=1.920064199e+00 la0=1.303350368e-07 wa0=-2.992883941e-07 pa0=-1.622753272e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-4.184869698e-01 lags=1.572962975e-06 wags=1.671892643e-06 pags=-3.909980840e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='5.608775762e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.581215293e-07 wvoff=-3.223580654e-07 pvoff=2.833651411e-13 nfactor='1.517998730e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.127144829e-06 wnfactor=2.343067921e-06 pnfactor=-2.071389050e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-7.195305916e-03 lpdiblc2=2.873909442e-08 wpdiblc2=2.784291210e-08 ppdiblc2=-6.056252642e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-1.454495035e-02 ldelta=6.084054077e-08 wdelta=2.069701677e-07 pdelta=-2.651730373e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.957152440e-01 lkt1=-2.788106283e-07 wkt1=-6.891615116e-07 pkt1=1.365068509e-12 kt2=9.507727976e-02 lkt2=-2.942021378e-07 wkt2=-4.577825797e-07 pkt2=8.971394105e-13 at=1.100532716e+06 lat=-1.649471019e+00 wat=-2.431414080e+00 pat=4.652861783e-6 ute=-0.13298 ua1=9.067491425e-10 lua1=-4.128392545e-16 wua1=-6.423835679e-16 pua1=1.258911197e-21 ub1=-9.396030676e-19 lub1=1.602532782e-24 wub1=2.493563087e-24 pub1=-4.886760259e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.21 pmos lmin=1e-06 lmax=1.5e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.171226900e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.078214540e-07 wvth0=-5.875180606e-08 pvth0=1.138138479e-13 k1=0.64774 k2=1.188401021e-01 lk2=-1.500605456e-07 wk2=-5.343008381e-07 pk2=6.960851484e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-2.903544755e+05 lvsat=4.085198429e-01 wvsat=1.262799853e+00 pvsat=-1.245739592e-6 ua=-3.166649539e-09 lua=-1.728755708e-16 wua=2.230295818e-16 pua=1.438852095e-21 ub=3.637729034e-18 lub=-1.542261147e-25 wub=-2.474351625e-24 pub=7.787490349e-31 uc=1.588070197e-10 luc=-9.127425744e-17 wuc=-5.194283692e-16 puc=5.574850778e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.956838409e-03 lu0=-1.051311271e-09 wu0=-5.691951688e-09 pu0=8.966831339e-15 a0=2.409537553e+00 la0=-5.841736916e-07 wa0=-1.555614159e-06 pa0=2.111682632e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=9.467218723e-01 lags=-4.199006327e-07 wags=-2.090488381e-06 pags=1.582154861e-12 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='1.501229882e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.981616283e-07 wvoff=-5.546870569e-07 pvoff=6.225073864e-13 nfactor='5.496423753e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-4.680361098e-06 wnfactor=-1.635256492e-05 pnfactor=2.521956099e-11 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.406441466e-02 lpdiblc2=3.876627591e-08 wpdiblc2=4.281495479e-08 ppdiblc2=-8.241796572e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.790876938e-02 ldelta=-1.572877660e-08 wdelta=-1.266175852e-07 pdelta=2.217816850e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.219204103e+00 lkt1=4.853522329e-07 wkt1=2.260496256e-06 pkt1=-2.940694416e-12 kt2=-2.421483668e-01 lkt2=1.980629998e-07 wkt2=4.577825797e-07 pkt2=-4.393568308e-13 at=-6.358975664e+05 lat=8.852830864e-01 wat=2.795073820e+00 pat=-2.976503929e-6 ute=-6.632089890e-01 lute=7.740017667e-07 wute=3.038182250e-06 pute=-4.434986540e-12 ua1=5.903123375e-10 lua1=4.907937160e-17 wua1=6.423835679e-16 pua1=-6.165276293e-22 ub1=4.828937376e-19 lub1=-4.739569296e-25 wub1=-2.493563087e-24 pub1=2.393197173e-30 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.22 pmos lmin=5e-07 lmax=1e-06 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.401848364e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.028744100e-08 wvth0=4.014122895e-08 pvth0=1.890125752e-14 k1=0.64774 k2=-6.016100630e-02 lk2=2.173576815e-08 wk2=3.663957825e-07 pk2=-1.683584333e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=3.764505238e+04 lvsat=9.372229596e-02 wvsat=3.172331587e-01 pvsat=-3.382319565e-7 ua=-3.837572347e-09 lua=4.710425946e-16 wua=3.302977849e-15 pua=-1.517128254e-21 ub=3.978470502e-18 lub=-4.812527382e-25 wub=-3.192019875e-24 pub=1.467531137e-30 uc=7.364656971e-11 luc=-9.541515599e-18 wuc=8.464167158e-17 puc=-2.227114383e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=7.950743415e-04 lu0=1.023441792e-09 wu0=7.557579452e-09 pu0=-3.749406173e-15 a0=1.585132203e+00 la0=2.070493436e-07 wa0=-1.311960025e-06 pa0=-2.267879137e-14 keta=-0.01258 a1=0.0 a2=0.46703705 ags=6.151373390e-01 lags=-1.016623768e-07 wags=-6.013236127e-07 pags=1.529289739e-13 b0=-1.318902119e-06 lb0=1.265816309e-12 wb0=4.614129815e-12 pb0=-4.428411089e-18 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.854608085e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-5.757563522e-09 wvoff=2.075048648e-07 pvoff=-1.090063105e-13 nfactor='7.515410873e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.264599603e-07 wnfactor=9.115829318e-06 pnfactor=7.762696187e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-7.163536690e-03 lpdiblc2=3.214315827e-08 wpdiblc2=-2.894381490e-08 ppdiblc2=-1.354748652e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.747194670e-03 ldelta=1.705779472e-08 wdelta=1.288737721e-07 pdelta=-2.342614519e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-4.739352872e-01 lkt1=-2.299195126e-07 wkt1=-6.344063283e-07 pkt1=-1.623116614e-13 kt2=-1.010471396e-02 lkt2=-2.464089603e-08 wkt2=-3.568552991e-08 pkt2=3.424918733e-14 at=5.003923223e+05 lat=-2.052711343e-01 wat=-6.130651057e-01 pat=2.944574051e-7 ute=5.911019272e-01 lute=-4.298231351e-07 wute=-2.784327241e-06 pute=1.153166944e-12 ua1=4.070694500e-10 lua1=2.249467329e-16 ub1=4.795829717e-19 lub1=-4.707794221e-25 wub1=2.544921246e-25 pub1=-2.442488166e-31 uc1=-2.194613080e-11 luc1=1.150272929e-17 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.23 pmos lmin=3.5e-07 lmax=5e-07 wmin=3.0e-06 wmax=5.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.003867407e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-5.398473349e-08 wvth0=-1.013581638e-06 pvth0=5.033503458e-13 k1=0.64774 k2=-1.020604929e-02 lk2=-1.231023330e-09 wk2=-3.996198136e-07 pk2=1.838172370e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=8.242000534e+05 lvsat=-2.678963658e-01 wvsat=-2.799214680e+00 pvsat=1.094554937e-6 ua=-2.881034865e-09 lua=3.127448699e-17 wua=1.092095741e-15 pua=-5.006752053e-22 ub=2.752719524e-18 lub=8.228627404e-26 wub=-1.497596022e-24 pub=6.885197713e-31 uc=-8.003748206e-12 luc=2.799721806e-17 wuc=3.116175797e-16 puc=-1.266233176e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.346949993e-03 lu0=3.099669611e-10 wu0=5.103780807e-09 pu0=-2.621272246e-15 a0=5.729119855e+00 la0=-1.698148980e-06 wa0=-1.202598461e-05 pa0=4.903094012e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-6.795654428e-02 lags=2.123900360e-07 wags=1.140037398e-06 pags=-6.476617509e-13 b0=4.396340397e-06 lb0=-1.361766438e-12 wb0=-1.538043272e-11 pb0=4.764089033e-18 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='6.980523652e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.119527451e-07 wvoff=-9.070632611e-08 pvoff=2.809628451e-14 nfactor='-1.580557337e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.485673410e-06 wnfactor=1.042545505e-05 pnfactor=1.741691893e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-2.097044619e-02 lpdiblc2=3.849088492e-08 wpdiblc2=-1.440059720e-07 ppdiblc2=3.935234022e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.786927005e-02 ldelta=-7.824829430e-09 wdelta=-1.077854093e-07 pdelta=8.537791347e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.437578448e+00 lkt1=2.131154305e-07 wkt1=1.535531919e-07 pkt1=-5.245760508e-13 kt2=-7.957261347e-02 lkt2=7.296970774e-09 wkt2=1.189517664e-07 pkt2=-3.684530963e-14 at=1.131592643e+05 lat=-2.724073588e-02 wat=8.400481814e-02 pat=-2.602049242e-8 ute=-2.308989607e-01 lute=-5.190822693e-08 wute=-8.461833648e-07 pute=2.621052972e-13 ua1=8.9635e-10 ub1=-4.312183725e-19 lub1=-5.203850413e-26 wub1=-8.483070821e-25 pub1=2.627631187e-31 uc1=3.0734e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.24 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.105726804e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=4.422444448e-8 k1=0.64774 k2=-1.043760653e-02 wk2=2.747387613e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.844218308e-09 wua=-4.416044384e-17 ub=2.872303364e-18 wub=7.104071401e-26 uc=5.901170046e-11 wuc=5.849658793e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.487440351e-03 wu0=-6.059260900e-11 a0=1.887787647e+00 wa0=-3.992200124e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.487466007e-01 wags=-2.640522539e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.650507143e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-5.315965429e-8 nfactor='2.594537465e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=5.389974173e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.696427525e-03 wpdiblc2=-1.368653756e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.473866424e-02 wdelta=-1.241612479e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.767537323e-01 wkt1=-1.620336285e-7 kt2=-0.055045 at=2.871894475e+05 wat=-1.356813637e-2 ute=-0.29175 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.25 pmos lmin=8e-06 lmax=2.0e-05 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.105726804e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=4.422444448e-8 k1=0.64774 k2=-1.043760653e-02 wk2=2.747387613e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.844218308e-09 wua=-4.416044384e-17 ub=2.872303364e-18 wub=7.104071401e-26 uc=5.901170046e-11 wuc=5.849658793e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.487440351e-03 wu0=-6.059260900e-11 a0=1.887787647e+00 wa0=-3.992200124e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.487466007e-01 wags=-2.640522539e-7 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.650507143e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-5.315965429e-8 nfactor='2.594537465e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=5.389974173e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.696427525e-03 wpdiblc2=-1.368653756e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.473866424e-02 wdelta=-1.241612479e-8 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.767537323e-01 wkt1=-1.620336285e-7 kt2=-0.055045 at=2.871894475e+05 wat=-1.356813637e-2 ute=-0.29175 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.26 pmos lmin=4e-06 lmax=8e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.496937149e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=3.113936547e-07 wvth0=8.005262258e-08 pvth0=-2.851833406e-13 k1=0.64774 k2=-2.898800927e-02 lk2=1.476565683e-07 wk2=5.318716717e-08 pk2=-2.046713683e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.824908567e-09 lua=-1.537007083e-16 wua=-1.248212545e-17 pua=-2.521514948e-22 ub=2.915415159e-18 lub=-3.431591099e-25 wub=-6.042430730e-26 pub=1.046428703e-30 uc=5.901170046e-11 wuc=5.849658793e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.668192565e-03 lu0=-1.438742434e-09 wu0=-2.683390210e-10 pu0=1.653609503e-15 a0=1.836740189e+00 la0=4.063250106e-07 wa0=-4.223483527e-07 pa0=1.840958063e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.412045154e-01 lags=6.003311312e-08 wags=-3.096959589e-07 pags=3.633124813e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.002264042e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=2.799896977e-07 wvoff=1.022636413e-08 pvoff=-5.045368601e-13 nfactor='2.743135622e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.182804182e-06 wnfactor=-2.343349416e-07 pnfactor=2.294276021e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.864751278e-03 lpdiblc2=-1.339814998e-09 wpdiblc2=-4.856278219e-09 ppdiblc2=2.776061882e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.940244608e-02 ldelta=4.247496246e-08 wdelta=-1.693978866e-08 pdelta=3.600723346e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-9.301727636e-01 lkt1=4.252021348e-07 wkt1=-2.542492134e-07 pkt1=7.340130013e-13 kt2=-0.055045 at=3.022161518e+05 lat=-1.196088098e-01 wat=-2.699974336e-02 pat=1.069122338e-7 ute=-4.489223769e-01 lute=1.251052827e-6 ua1=6.683900700e-10 lua1=1.096847978e-16 ub1=-1.521398367e-19 lub1=1.599779781e-26 wub1=-7.914986241e-26 pub1=6.300131173e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.27 pmos lmin=2e-06 lmax=4e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.910634709e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=7.923254614e-08 wvth0=3.567267253e-08 pvth0=-1.094498334e-13 k1=0.64774 k2=9.756400293e-03 lk2=-5.761607532e-09 wk2=3.725513444e-09 pk2=-8.815584993e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.838017356e-09 lua=-1.017931809e-16 wua=-1.545515533e-16 pua=3.104079223e-22 ub=2.797647912e-18 lub=1.231697489e-25 wub=2.986949021e-25 pub=-3.755935860e-31 uc=7.357684716e-11 luc=-5.767433966e-17 wuc=-9.434977028e-18 puc=6.052333669e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.390816923e-03 lu0=-3.404042337e-10 wu0=-3.333800107e-11 pu0=7.230642142e-16 a0=2.187557701e+00 la0=-9.828246334e-07 wa0=-5.374623224e-07 pa0=6.399183481e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=4.113887699e-01 lags=-2.178789884e-07 wags=-3.655607153e-07 pags=5.845229503e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.534680530e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=9.483831656e-08 wvoff=-1.458347556e-07 pvoff=1.134261589e-13 nfactor='2.442390998e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=8.069342165e-09 wnfactor=4.788224695e-07 pnfactor=-5.296490378e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=5.084365503e-05 lpdiblc2=9.802555713e-09 wpdiblc2=4.335773577e-11 ppdiblc2=8.359285348e-15 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.225946006e-02 ldelta=7.075940138e-08 wdelta=9.462207101e-09 pdelta=-6.853806924e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.359719254e-01 lkt1=5.219036575e-08 wkt1=-5.803140725e-08 pkt1=-4.296045645e-14 kt2=-0.055045 at=3.032778113e+05 lat=-1.238127156e-1 ute=-1.439208871e-01 lute=4.332317780e-08 wute=3.336311932e-08 pute=-1.321096117e-13 ua1=6.9609e-10 ub1=-1.737917953e-19 lub1=1.017341409e-25 wub1=1.582997248e-25 pub1=-3.102278857e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.28 pmos lmin=1.5e-06 lmax=2e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-1.285149702e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-2.393218782e-07 wvth0=-1.483271916e-07 pvth0=2.511439003e-13 k1=0.64774 k2=4.848559869e-02 lk2=-8.166115410e-08 wk2=-4.450035046e-08 pk2=8.569505179e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.889959278e-09 wua=3.840038595e-18 ub=2.860497637e-18 wub=1.070410758e-25 uc=4.414740990e-11 wuc=2.144821557e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.962145310e-03 lu0=4.996849596e-10 wu0=6.031883984e-10 pu0=-5.243683972e-16 a0=1.998671518e+00 la0=-6.126549356e-07 wa0=-5.389933932e-07 pa0=6.429188641e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=7.400714333e-02 lags=4.433046542e-07 wags=1.700820798e-07 pags=-4.652030175e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='2.344909640e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-2.518750670e-07 wvoff=-2.228297972e-07 pvoff=2.643171916e-13 nfactor='2.098065076e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=6.828620682e-07 wnfactor=5.742147648e-07 pnfactor=-7.165940886e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.854832885e-03 lpdiblc2=1.353720531e-08 wpdiblc2=1.155768432e-08 ppdiblc2=-1.420591618e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=6.868625346e-02 ldelta=-3.982300699e-08 wdelta=-4.683489872e-08 pdelta=4.179018389e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-9.407003871e-01 lkt1=2.574319685e-07 wkt1=5.789569389e-08 pkt1=-2.701485929e-13 kt2=-0.055045 at=3.362938622e+05 lat=-1.885159214e-01 wat=-1.009456466e-01 pat=1.978282309e-7 ute=-1.218144053e-01 wute=-3.404834221e-8 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.29 pmos lmin=1e-06 lmax=1.5e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-1.583172225e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-1.958180403e-07 wvth0=-2.380730808e-07 pvth0=3.821504621e-13 k1=0.64774 k2=-6.095782474e-02 lk2=7.809888326e-08 wk2=1.397460045e-08 pk2=3.362421945e-16 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.202233871e-09 lua=4.558428375e-16 wua=3.315403722e-16 pua=-4.783605620e-22 ub=2.754845221e-18 lub=1.542261147e-25 wub=2.179125102e-25 pub=-1.618445763e-31 uc=-5.146949015e-11 luc=1.395767699e-16 wuc=1.217883993e-16 puc=-1.464715831e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.543667671e-04 lu0=2.992614687e-09 wu0=2.548959931e-09 pu0=-3.364708391e-15 a0=2.089856574e+00 la0=-7.457623219e-07 wa0=-5.807796204e-07 pa0=7.039163092e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=2.438070685e-01 lags=1.954392135e-07 wags=5.297861567e-08 pags=-2.942612357e-13 b0=0.0 b1=2.1073e-24 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-8.465912969e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-9.406408397e-08 wvoff=-2.507492022e-07 pvoff=3.050725430e-13 nfactor='-1.442187161e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=5.850745271e-06 wnfactor=4.806021324e-06 pnfactor=-6.893973713e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=3.828704778e-03 lpdiblc2=5.240661209e-09 wpdiblc2=-1.174828784e-08 ppdiblc2=1.981497668e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=4.732044066e-03 ldelta=5.353415017e-08 wdelta=-2.544854537e-08 pdelta=1.057145459e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-2.341822281e-01 lkt1=-7.739079140e-07 wkt1=-7.432274779e-07 pkt1=8.992909571e-13 kt2=-9.202608700e-02 lkt2=5.398314175e-8 at=2.257723765e+05 lat=-2.718218264e-02 wat=1.674992195e-01 pat=-1.940341623e-7 ute=5.842142473e-01 lute=-1.030625326e-06 wute=-7.657076719e-07 pute=1.068039706e-12 ua1=8.009714800e-10 lua1=-1.531007404e-16 ub1=-3.348293300e-19 lub1=3.108527845e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.30 pmos lmin=5e-07 lmax=1e-06 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.545819229e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=-7.452994104e-09 wvth0=8.404367589e-08 pvth0=7.299890484e-14 k1=0.64774 k2=7.088170267e-02 lk2=-4.843410317e-08 wk2=-3.320559214e-08 pk2=4.561743203e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.354232840e+05 lvsat=-1.119383679e-02 wvsat=1.906841485e-02 pvsat=-1.830091115e-8 ua=-2.704513502e-09 lua=-2.184428689e-17 wua=-1.521695294e-16 pua=-1.411998392e-23 ub=2.954136129e-18 lub=-3.704333489e-26 wub=-6.841668763e-26 pub=1.129598713e-31 uc=1.169824067e-10 luc=-2.209493814e-17 wuc=-4.750654307e-17 puc=1.600923776e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.612409315e-03 lu0=-2.302666479e-10 wu0=-1.033596180e-09 pu0=7.364983610e-17 a0=8.530955995e-01 la0=4.412190234e-07 wa0=9.203109281e-07 pa0=-7.367553447e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=5.539794167e-01 lags=-1.022486978e-07 wags=-4.148287669e-07 pags=1.547168998e-13 b0=5.068653630e-07 lb0=-4.864640321e-13 wb0=-9.533618939e-13 pb0=9.149890777e-19 b1=2.325991428e-07 lb1=-2.232370273e-13 wb1=-7.092873608e-13 pb1=6.807385445e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.079762787e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-7.168545017e-08 wvoff=-2.877630522e-08 pvoff=9.203405516e-14 nfactor='4.134546827e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=4.984748262e-07 wnfactor=-1.200301618e-06 pnfactor=-1.129405269e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.938584188e-02 lpdiblc2=2.752082236e-08 wpdiblc2=8.326858090e-09 ppdiblc2=5.478553759e-16 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=5.288997439e-02 ldelta=7.314576543e-09 wdelta=-2.098212208e-08 pdelta=6.284804841e-15 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.404588832e-01 lkt1=-2.880088943e-07 wkt1=1.783301923e-07 pkt1=1.482598311e-14 kt2=-2.180719750e-02 lkt2=-1.340943745e-8 at=3.201167328e+05 lat=-1.177291786e-01 wat=-6.333308374e-02 pat=2.750714066e-8 ute=-4.440801196e-01 lute=-4.371980700e-08 wute=3.723548224e-07 pute=-2.421577241e-14 ua1=4.070694500e-10 lua1=2.249467329e-16 ub1=5.630394850e-19 lub1=-5.508768107e-25 wub1=-2.869859255e-41 pub1=2.736911063e-47 uc1=-2.194613080e-11 luc1=1.150272929e-17 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.31 pmos lmin=3.5e-07 lmax=5e-07 wmin=1e-06 wmax=3.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-6.407084496e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' lvth0=1.240936765e-07 wvth0=3.291345000e-07 pvth0=-3.968160155e-14 k1=0.64774 k2=-1.531870269e-01 lk2=5.458149526e-08 wk2=3.638609370e-08 pk2=1.362265447e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-1.398632840e+05 lvsat=1.153691628e-01 wvsat=1.405981331e-01 pvsat=-7.417419912e-8 ua=-2.354576561e-09 lua=-1.827277954e-16 wua=-5.132851588e-16 pua=1.519029267e-22 ub=2.093061851e-18 lub=3.588355646e-25 wub=5.139627657e-25 pub=-1.547890823e-31 uc=1.137836906e-10 luc=-2.062432842e-17 wuc=-5.976079263e-17 puc=2.164312900e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=4.588194344e-03 lu0=-6.788838153e-10 wu0=-1.730665234e-09 pu0=3.941273337e-16 a0=2.112123481e+00 la0=-1.376190449e-07 wa0=-9.963231017e-07 pa0=1.444171505e-13 keta=-1.176195491e-02 lketa=-3.760962317e-10 wketa=-2.494545072e-09 pketa=1.146867097e-15 a1=0.0 a2=0.46703705 ags=3.315787691e-01 wags=-7.830478701e-8 b0=-1.642697271e-06 lb0=5.017973888e-13 wb0=3.034996672e-12 pb0=-9.186587729e-19 b1=-5.551192378e-07 lb1=1.389164982e-13 wb1=1.692779494e-12 pb1=-4.236116918e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='4.960232045e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.493742126e-07 wvoff=5.253609922e-07 pvoff=-1.627305673e-13 nfactor='-1.025751707e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=7.115226203e-06 wnfactor=-6.492776729e-06 pnfactor=1.303810163e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-8.380581845e-02 lpdiblc2=5.713790659e-08 wpdiblc2=4.760408645e-08 ppdiblc2=-1.750985036e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-8.821774543e-03 ldelta=3.568655312e-08 wdelta=9.558212866e-08 pdelta=-4.730560944e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.483864833e+00 lkt1=5.377199103e-08 wkt1=2.946988019e-07 pkt1=-3.867448514e-14 kt2=-7.233698973e-02 lkt2=9.821634527e-09 wkt2=9.688746978e-08 pkt2=-4.454401423e-14 at=1.424300879e+05 lat=-3.603774366e-02 wat=-5.253572802e-03 pat=8.050855116e-10 ute=-6.280372522e-01 lute=4.085448470e-08 wute=3.648493470e-07 pute=-2.076513008e-14 ua1=7.087088751e-10 lua1=8.626800716e-17 wua1=5.721924709e-16 pua1=-2.630654885e-22 ub1=-3.120318652e-19 lub1=-1.485627575e-25 wub1=-1.211754179e-24 pub1=5.571039838e-31 uc1=3.224846359e-11 luc1=-1.341323549e-17 wuc1=-8.896638057e-17 puc1=4.090229347e-23 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.32 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.885964127e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))' wvth0=2.116259317e-8 k1=0.64774 k2=1.799007650e-02 wk2=-2.358077587e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.694093041e-09 wua=-2.017015980e-16 ub=2.757516609e-18 wub=1.914977057e-25 uc=7.060795191e-11 wuc=-6.319424287e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.968132563e-03 wu0=-5.650300552e-10 a0=1.218929682e+00 wa0=3.026781984e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-1.259666076e-01 wags=2.341108375e-7 b0=-2.149574428e-07 wb0=2.255759105e-13 b1=-2.238818130e-07 wb1=2.349411268e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.757161654e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-4.196735120e-8 nfactor='2.712795481e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=-7.019998375e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.669956697e-03 wpdiblc2=-1.340875322e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.201855896e-02 wdelta=9.323282458e-10 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.128568835e+00 wkt1=1.022206366e-7 kt2=-0.055045 at=2.636706353e+05 wat=1.111245810e-2 ute=-2.995155341e-01 wute=8.149135942e-9 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.33 pmos lmin=8e-06 lmax=2.0e-05 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.885964127e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=2.116259317e-8 k1=0.64774 k2=1.799007650e-02 wk2=-2.358077587e-9 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.694093041e-09 wua=-2.017015980e-16 ub=2.757516609e-18 wub=1.914977057e-25 uc=7.060795191e-11 wuc=-6.319424287e-18 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.968132563e-03 wu0=-5.650300552e-10 a0=1.218929682e+00 wa0=3.026781984e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-1.259666076e-01 wags=2.341108375e-7 b0=-2.149574428e-07 wb0=2.255759105e-13 b1=-2.238818130e-07 wb1=2.349411268e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.757161654e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-4.196735120e-8 nfactor='2.712795481e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=-7.019998375e-8 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=2.669956697e-03 wpdiblc2=-1.340875322e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.201855896e-02 wdelta=9.323282458e-10 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.128568835e+00 wkt1=1.022206366e-7 kt2=-0.055045 at=2.636706353e+05 wat=1.111245810e-2 ute=-2.995155341e-01 wute=8.149135942e-9 ua1=6.8217e-10 ub1=-1.5013e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.34 pmos lmin=4e-06 lmax=8e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.442736304e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-3.527982668e-07 wvth0=-3.057500330e-08 pvth0=4.118183335e-13 k1=0.64774 k2=5.616896773e-02 lk2=-3.038944295e-07 wk2=-3.617639419e-08 pk2=2.691853456e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.631805821e-09 lua=-4.957907057e-16 wua=-2.151237613e-16 pua=1.068370643e-22 ub=2.606521276e-18 lub=1.201885103e-24 wub=2.637283164e-25 pub=-5.749376039e-31 uc=6.347964166e-11 luc=5.673956748e-17 wuc=1.161010228e-18 puc=-5.954238863e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.822447098e-03 lu0=1.159619887e-09 wu0=-4.302134191e-10 pu0=-1.073106719e-15 a0=1.002999487e+00 la0=1.718750369e-06 wa0=4.525774716e-07 pa0=-1.193160740e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-2.798751262e-01 lags=1.225073331e-06 wags=3.420637748e-07 pags=-8.592783928e-13 b0=-1.103930694e-07 lb0=-8.323062710e-13 wb0=1.158462662e-13 pb0=8.734205362e-19 b1=-1.162055617e-07 lb1=-8.570760415e-13 wb1=1.219458840e-13 pb1=8.994138838e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.344037361e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.291674734e-06 wvoff=-1.857865228e-07 pvoff=1.144764651e-12 nfactor='2.378145409e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.663730907e-06 wnfactor=1.486850576e-07 pnfactor=-1.742270208e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=-1.201194122e-03 lpdiblc2=3.081339272e-08 wpdiblc2=-5.894832481e-10 ppdiblc2=-5.980893059e-15 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-4.572089290e-03 ldelta=1.320574124e-07 wdelta=8.219040816e-09 pdelta=-5.800041038e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.349241874e+00 lkt1=1.756502221e-06 wkt1=1.855210728e-07 pkt1=-6.630506466e-13 kt2=-0.055045 at=2.517890566e+05 lat=9.457439664e-02 wat=2.591834958e-02 pat=-1.178511947e-7 ute=-4.152788368e-01 lute=9.214469487e-07 wute=-3.530546367e-08 pute=3.458877493e-13 ua1=6.683900700e-10 lua1=1.096847978e-16 ub1=-2.934552795e-19 lub1=1.140833394e-24 wub1=6.914628064e-26 pub1=-5.503871073e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.35 pmos lmin=2e-06 lmax=4e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.026457489e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-1.216592704e-07 wvth0=4.782709189e-08 pvth0=1.013656371e-13 k1=0.64774 k2=-1.879107063e-02 lk2=-7.071417546e-09 wk2=3.368317234e-08 pk2=-7.441072983e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.884318497e-09 lua=5.040963646e-16 wua=-1.059632286e-16 pua=-3.254113550e-22 ub=3.074396941e-18 lub=-6.507855606e-25 wub=8.275024716e-27 pub=4.365935679e-31 uc=7.780871988e-11 wuc=-1.387589580e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.943398719e-03 lu0=6.806817034e-10 wu0=-6.132162332e-10 pu0=-3.484613259e-16 a0=1.656740828e+00 la0=-8.699019034e-07 wa0=1.957584248e-08 pa0=5.214174611e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=-6.453393875e-02 lags=3.723760636e-07 wags=1.338716232e-07 pags=-3.488952077e-14 b0=-3.773082106e-07 lb0=2.246109593e-13 wb0=3.959464815e-13 pb0=-2.357062914e-19 b1=-3.511601521e-07 lb1=7.328539813e-14 wb1=3.685067613e-13 pb1=-7.690555022e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-4.344406320e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=3.753810393e-07 wvoff=1.490173069e-07 pvoff=-1.809748133e-13 nfactor='3.258141797e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-8.208347904e-07 wnfactor=-3.772247875e-07 pnfactor=3.402013010e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.447540278e-03 lpdiblc2=2.032506669e-08 wpdiblc2=-1.422332907e-09 ppdiblc2=-2.683016622e-15 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.405204175e-02 ldelta=-2.088449046e-08 wdelta=-1.340688454e-08 pdelta=2.763284756e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.381838008e-01 lkt1=-2.671599837e-07 wkt1=-5.571026967e-08 pkt1=2.921651615e-13 kt2=-0.055045 at=3.001146598e+05 lat=-9.678291079e-02 wat=3.319404806e-03 pat=-2.836502311e-8 ute=-1.339493575e-01 lute=-1.925474569e-07 wute=2.289901608e-08 pute=1.154125606e-13 ua1=6.9609e-10 ub1=1.088390903e-19 lub1=-4.521517372e-25 wub1=-1.382925613e-25 pub1=2.710188470e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.36 pmos lmin=1.5e-06 lmax=2e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.647247235e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=9.955085108e-8 k1=0.64774 k2=-2.239939697e-02 wk2=2.988622223e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-2.627093665e-09 wua=-2.720106097e-16 ub=2.742321135e-18 wub=2.310552609e-25 uc=7.780871988e-11 wuc=-1.387589580e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.290729605e-03 wu0=-7.910253037e-10 a0=1.212856708e+00 wa0=2.856390960e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=1.254780851e-01 wags=1.160685765e-7 b0=-2.626961635e-07 wb0=2.756728285e-13 b1=-3.137648731e-07 wb1=3.292642303e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-2.428952618e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=5.667143963e-8 nfactor='2.839295113e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=-2.036305530e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.181879512e-02 wpdiblc2=-2.791393564e-9 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.339533020e-02 wdelta=6.933055621e-10 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-9.745073031e-01 wkt1=9.337260393e-8 kt2=-0.055045 at=2.507293245e+05 wat=-1.115439191e-2 ute=-2.322003879e-01 wute=8.179048722e-8 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.37 pmos lmin=1e-06 lmax=1.5e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-6.396671517e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=4.013472096e-07 wvth0=2.670545722e-07 pvth0=-2.445135568e-13 k1=0.64774 k2=-1.203013508e-01 lk2=1.429123771e-07 wk2=7.624957799e-08 pk2=-6.767890857e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=4.632068748e+04 lvsat=1.130420365e-01 wvsat=8.126465968e-02 pvsat=-1.186260870e-7 ua=-1.827593103e-09 lua=-1.167070946e-15 wua=-1.111004901e-15 pua=1.224721916e-21 ub=1.881969554e-18 lub=1.255898219e-24 wub=1.133906489e-24 pub=-1.317937080e-30 uc=1.248148530e-10 luc=-6.861720286e-17 wuc=-6.320403791e-17 puc=7.200675545e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=5.307352675e-03 lu0=-2.943765527e-09 wu0=-2.753633375e-09 pu0=2.864917132e-15 a0=3.843372598e-01 la0=1.209431265e-06 wa0=1.208988937e-06 pa0=-1.347859930e-12 keta=-1.064964207e-02 lketa=-2.817839987e-09 wketa=-2.025713750e-09 pketa=2.957035647e-15 a1=0.0 a2=0.46703705 ags=6.469856093e-01 lags=-7.612706086e-07 wags=-3.701161388e-07 pags=7.097081382e-13 b0=9.270702054e-08 lb0=-5.187997978e-13 wb0=-9.728656194e-14 pb0=5.444274703e-19 b1=-7.387666930e-09 lb1=-4.472341267e-13 wb1=7.752602901e-15 pb1=4.693265980e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-5.093191458e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=3.889122647e-07 wvoff=1.948881694e-07 pvoff=-2.017618713e-13 nfactor='4.025305005e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.731277940e-06 wnfactor=-9.315540199e-07 pnfactor=1.062586281e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=6.589225566e-03 lpdiblc2=7.633864163e-09 wpdiblc2=-1.464517283e-08 ppdiblc2=1.730355429e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-6.080112907e-02 ldelta=1.229057814e-07 wdelta=4.332183544e-08 pdelta=-6.222699649e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.114035943e+00 lkt1=2.036769322e-07 wkt1=1.800892508e-07 pkt1=-1.265846253e-13 kt2=-2.187393836e-01 lkt2=2.389528765e-07 wkt2=1.329726801e-07 pkt2=-1.941068697e-13 at=2.789164211e+05 lat=-4.114611415e-02 wat=1.117299654e-01 pat=-1.793804405e-7 ute=-2.225308097e-01 lute=-1.411516677e-08 wute=8.088897753e-08 pute=1.315978778e-15 ua1=1.009910354e-09 lua1=-4.580992619e-16 wua1=-2.192600366e-16 pua1=3.200648385e-22 ub1=-5.470613180e-19 lub1=6.206584290e-25 wub1=2.227158238e-25 pub1=-3.251094238e-31 uc1=9.220990490e-11 luc1=-1.491439784e-16 wuc1=-1.072179433e-16 puc1=1.565113927e-22 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.38 pmos lmin=5e-07 lmax=1e-06 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.520389329e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=1.252960266e-07 wvth0=8.137506719e-08 pvth0=-6.630765196e-14 k1=0.64774 k2=3.039875831e-02 lk2=-1.722052628e-09 wk2=9.277128716e-09 pk2=-3.402100385e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=2.024570779e+05 lvsat=-3.680986426e-02 wvsat=-5.127671443e-02 pvsat=8.580496838e-9 ua=-3.126366219e-09 lua=7.942655241e-17 wua=2.905218682e-16 pua=-1.203934001e-22 ub=3.371974735e-18 lub=-1.741342528e-25 wub=-5.068956849e-25 pub=2.568228064e-31 uc=6.331084342e-11 luc=-9.588729639e-18 wuc=8.816288089e-18 puc=2.885247571e-24 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.423904107e-03 lu0=-1.763757634e-10 wu0=2.136188077e-10 pu0=1.709684965e-17 a0=2.087495250e+00 la0=-4.251746161e-07 wa0=-3.750655962e-07 pa0=1.724364078e-13 keta=-1.358565664e-02 wketa=1.055334071e-9 a1=0.0 a2=0.46703705 ags=-2.192589803e-01 lags=7.010763632e-08 wags=3.966060604e-07 pags=-2.615349252e-14 b0=-1.503845609e-06 lb0=1.013491588e-12 wb0=1.156674178e-12 pb0=-6.590613503e-19 b1=-1.473164503e-06 lb1=9.595451921e-13 wb1=1.080737598e-12 pb1=-5.604707509e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.440859299e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=3.837968566e-08 wvoff=9.117090449e-09 pvoff=-2.346807825e-14 nfactor='3.463380473e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.191970871e-06 wnfactor=-4.959809887e-07 pnfactor=6.445450641e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=1.609295702e-02 lpdiblc2=-1.487342103e-09 wpdiblc2=-2.890452252e-08 ppdiblc2=3.098896515e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=3.875671355e-02 ldelta=2.735514197e-08 wdelta=-6.150706422e-09 pdelta=-1.474572444e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-8.112745319e-01 lkt1=-8.689833222e-08 wkt1=2.526439924e-07 pkt1=-1.962190385e-13 kt2=6.281688107e-02 lkt2=-3.127074853e-08 wkt2=-8.880433880e-08 pkt2=1.874362413e-14 at=4.456865844e+05 lat=-2.012037784e-01 wat=-1.951058348e-01 pat=1.151052187e-7 ute=-7.493814870e-02 lute=-1.557672232e-07 wute=-1.502202354e-08 pute=9.336656205e-14 ua1=-1.397507771e-11 lua1=5.245747813e-16 wua1=4.418432853e-16 pua1=-3.144290747e-22 ub1=1.211546764e-18 lub1=-1.067165678e-24 wub1=-6.805422414e-25 pub1=5.417925043e-31 uc1=-9.113814615e-11 luc1=2.682431357e-17 wuc1=7.260996253e-17 puc1=-1.607843991e-23 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.39 pmos lmin=3.5e-07 lmax=5e-07 wmin=5.5e-07 wmax=1.0e-6 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-2.473877453e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=7.718264311e-08 wvth0=-8.361546036e-08 pvth0=9.546743084e-15 k1=0.64774 k2=-1.579111499e-01 lk2=8.485342766e-08 wk2=4.134357888e-08 pk2=-1.814465085e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=3.353436604e+04 lvsat=4.085235252e-02 wvsat=-4.136501404e-02 pvsat=4.023592582e-9 ua=-3.090501461e-09 lua=6.293772985e-17 wua=2.589929590e-16 pua=-1.058979842e-22 ub=2.660073422e-18 lub=1.531623757e-25 wub=-8.105804344e-26 pub=6.104395078e-32 uc=1.431885505e-11 luc=1.293533702e-17 wuc=4.461740688e-17 puc=-1.357431679e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.126749772e-03 lu0=-3.975905814e-11 wu0=8.523697766e-10 pu0=-2.765689083e-16 a0=1.1627 keta=-1.722141262e-02 lketa=1.671538808e-09 wketa=3.234598929e-09 pketa=-1.001917018e-15 a1=0.0 a2=0.46703705 ags=-7.847497015e-01 lags=3.300919954e-07 wags=1.093168077e-06 pags=-3.463978798e-13 b0=1.939084068e-06 lb0=-5.693953306e-13 wb0=-7.237175015e-13 pb0=2.054487245e-19 b1=9.030021305e-07 lb1=-1.328974178e-13 wb1=1.626298459e-13 pb1=-1.383707119e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='1.119114696e+00+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-5.423768021e-07 wvoff=-1.285099728e-07 pvoff=3.980596408e-14 nfactor='-1.909073582e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=9.177284096e-06 wnfactor=2.776785364e-06 pnfactor=-8.601092664e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=0.030097 pdiblc1=0.0 pdiblc2=3.792390015e-03 lpdiblc2=4.167843579e-09 wpdiblc2=-4.432129831e-08 ppdiblc2=3.807682782e-14 pdiblcb=-0.025 drout=0.43496 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.528726402e-01 ldelta=-2.510965531e-08 wdelta=-7.409966679e-08 pdelta=1.649381009e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.137205752e+00 lkt1=6.294854608e-08 wkt1=-6.908454456e-08 pkt1=-4.830434366e-14 kt2=1.602871186e-01 lkt2=-7.608269023e-08 wkt2=-1.472278042e-07 pkt2=4.560381236e-14 at=-5.965818746e+04 lat=3.112848044e-02 wat=2.068174592e-01 pat=-6.967901573e-8 ute=-8.296308305e-01 lute=1.912027372e-07 wute=5.764012449e-07 pute=-1.785402856e-13 ua1=1.960985545e-09 lua1=-3.834133652e-16 wua1=-7.419441622e-16 pua1=2.298172042e-22 ub1=-2.920996469e-18 lub1=8.327710739e-25 wub1=1.526088059e-24 pub1=-4.727057762e-31 uc1=-1.624596608e-10 luc1=5.961437994e-17 wuc1=1.153599358e-16 puc1=-3.573274011e-23 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.40 pmos lmin=2.0e-05 lmax=1.0e-04 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.041982960e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=-1.335879344e-7 k1=0.64774 k2=6.563561869e-02 wk2=-3.091672028e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.406118400e-09 wua=2.250849779e-16 ub=3.775680869e-18 wub=-4.187879157e-25 uc=5.984835477e-11 wuc=1.298567180e-19 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.511082007e-03 wu0=3.083231342e-10 a0=2.092557968e+00 wa0=-2.209728485e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=6.697004740e-01 wags=-2.428104199e-7 b0=8.358146572e-07 wb0=-4.042547846e-13 b1=-9.412157966e-07 wb1=6.649096819e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='4.228279606e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-4.007335033e-7 nfactor='-1.232836923e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=8.945444064e-6 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-5.291112804e-01 wpclm=3.351883249e-7 pdiblc1=0.0 pdiblc2=1.516110046e-03 wpdiblc2=-6.492619474e-10 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=9.797151477e-03 wdelta=2.263835451e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-7.406987260e-01 wkt1=-1.302679310e-7 kt2=-0.055045 at=2.535045069e+05 wat=1.720601514e-2 ute=-6.782284054e-01 wute=2.351488736e-7 ua1=6.8217e-10 ub1=-5.798356185e-20 wub1=-5.523239074e-26 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.41 pmos lmin=8e-06 lmax=2.0e-05 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='1.782232670e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-4.164464047e-06 wvth0=-2.586481892e-07 pvth0=2.496171421e-12 k1=0.64774 k2=1.244917779e-01 lk2=-1.174754224e-06 wk2=-6.619498442e-08 pk2=7.041453326e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.406118400e-09 wua=2.250849779e-16 ub=3.775680869e-18 wub=-4.187879157e-25 uc=5.984835477e-11 wuc=1.298567180e-19 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.324387223e-03 lu0=3.726381207e-09 wu0=4.202276141e-10 pu0=-2.233585443e-15 a0=1.688032644e+00 la0=8.074224322e-06 wa0=2.149882123e-08 pa0=-4.839673910e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=6.697004740e-01 wags=-2.428104199e-7 b0=1.156596772e-06 lb0=-6.402730815e-12 wb0=-5.965309426e-13 pb0=3.837784045e-18 b1=-2.039824185e-06 lb1=2.192794878e-11 wb1=1.323413353e-12 pb1=-1.314356864e-17 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='9.917979773e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-1.135649929e-05 wvoff=-7.417729933e-07 pvoff=6.807062961e-12 nfactor='-2.231374752e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=1.993056542e-04 wnfactor=1.493065984e-05 pnfactor=-1.194634105e-10 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-5.291112804e-01 wpclm=3.351883249e-7 pdiblc1=0.0 pdiblc2=4.126891095e-03 lpdiblc2=-5.211053704e-08 wpdiblc2=-2.214158887e-09 ppdiblc2=3.123495168e-14 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.316397107e-02 ldelta=-2.667983774e-07 wdelta=-5.748209480e-09 pdelta=1.599184138e-13 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-4.843556511e-01 lkt1=-5.116543690e-06 wkt1=-2.839194574e-07 pkt1=3.066846055e-12 kt2=-0.055045 at=2.141776519e+05 lat=7.849541940e-01 wat=4.077845337e-02 pat=-4.704999740e-7 ute=-6.782284054e-01 wute=2.351488736e-7 ua1=6.8217e-10 ub1=3.138322412e-21 lub1=-1.219977529e-24 wub1=-9.186872592e-26 pub1=7.312520911e-31 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.42 pmos lmin=4e-06 lmax=8e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-6.047853824e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=2.068089050e-06 wvth0=1.855150199e-07 pvth0=-1.039256682e-12 k1=0.64774 k2=-1.188872547e-01 lk2=7.624820310e-07 wk2=6.875195545e-08 pk2=-3.699985721e-13 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.472384212e-09 lua=5.274592941e-16 wua=2.887172452e-16 pua=-5.064969391e-22 ub=4.176623365e-18 lub=-3.191402030e-24 wub=-6.773877357e-25 pub=2.058389917e-30 uc=1.060162661e-10 luc=-3.674850325e-16 wuc=-2.433535741e-17 puc=1.947369881e-22 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=2.401861447e-03 lu0=-4.850044245e-09 wu0=-1.781152214e-10 pu0=2.529073942e-15 a0=3.101515483e+00 la0=-3.176745702e-06 wa0=-8.052688190e-07 pa0=1.741189814e-12 keta=-0.01258 a1=0.0 a2=0.46703705 ags=7.904733903e-01 lags=-9.613222203e-07 wags=-2.995009853e-07 pags=4.512427275e-13 b0=-1.802201028e-07 lb0=4.237997303e-12 wb0=1.577004504e-13 pb0=-2.165709286e-18 b1=9.534158330e-07 lb1=-1.897493456e-12 wb1=-5.191830407e-13 pb1=1.523038001e-18 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-7.704717858e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=2.670727457e-06 wvoff=2.679765916e-07 pvoff=-1.230291297e-12 nfactor='3.014385847e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-2.299955323e-06 wnfactor=-2.326761882e-07 pnfactor=1.232953391e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-5.291112804e-01 wpclm=3.351883249e-7 pdiblc1=0.0 pdiblc2=2.122913568e-03 lpdiblc2=-3.615937692e-08 wpdiblc2=-2.581946749e-09 ppdiblc2=3.416245112e-14 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-6.249104903e-03 ldelta=-3.267764591e-08 wdelta=9.224240621e-09 pdelta=4.074145412e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.151309080e+00 lkt1=1.922388645e-07 wkt1=6.688055187e-08 pkt1=2.745656808e-13 kt2=-0.055045 at=3.558881185e+05 lat=-3.430256922e-01 wat=-3.647841994e-02 pat=1.444454234e-7 ute=-1.254849582e+00 lute=4.589760407e-06 wute=4.679315616e-07 pute=-1.852892001e-12 ua1=6.683900700e-10 lua1=1.096847978e-16 ub1=-1.780957344e-19 lub1=2.226002542e-25 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.43 pmos lmin=2e-06 lmax=4e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-7.591661304e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-2.609905964e-08 wvth0=-8.807389870e-08 pvth0=4.408703787e-14 k1=0.64774 k2=8.549107185e-02 lk2=-4.680504776e-08 wk2=-2.882333530e-08 pk2=1.637518550e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.293999387e-09 lua=-1.789000171e-16 wua=1.395986772e-16 pua=8.397531024e-23 ub=3.280303632e-18 lub=3.578000342e-25 wub=-1.151450340e-25 pub=-1.679506205e-31 uc=1.321115660e-11 wuc=2.484375444e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.381987118e-03 lu0=-8.115968713e-10 wu0=3.226907574e-10 pu0=5.460074672e-16 a0=2.060081615e+00 la0=9.470720576e-07 wa0=-2.221858185e-07 pa0=-5.676730972e-13 keta=-0.01258 a1=0.0 a2=0.46703705 ags=3.760153667e-01 lags=6.798279386e-07 wags=-1.301927493e-07 pags=-2.191755597e-13 b0=1.250895750e-06 lb0=-1.428863693e-12 wb0=-5.799957158e-13 pb0=7.553831082e-19 b1=4.720168963e-07 lb1=8.725983406e-15 wb1=-1.249039152e-13 pb1=-3.820876616e-20 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.339007711e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=1.500653815e-07 wvoff=-3.112568474e-08 pvoff=-4.592105865e-14 nfactor='2.794417443e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=-1.428935434e-06 wnfactor=-9.926933684e-08 pnfactor=7.046956109e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-5.291112804e-01 wpclm=3.351883249e-7 pdiblc1=0.0 pdiblc2=-1.923241407e-02 lpdiblc2=4.840238170e-08 wpdiblc2=1.097319037e-08 ppdiblc2=-1.951250309e-14 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=-5.727314582e-02 ldelta=1.693648001e-07 wdelta=4.133325024e-08 pdelta=-8.640219670e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.528189248e+00 lkt1=1.684590112e-06 wkt1=3.578776157e-07 pkt1=-8.777099426e-13 kt2=-0.055045 at=3.056525575e+05 lat=-1.441054296e-1 ute=-1.499636517e-01 lute=2.146883463e-07 wute=3.249795199e-08 pute=-1.286837654e-13 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.44 pmos lmin=1.5e-06 lmax=2e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-8.923415846e-02+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' wvth0=-6.557764261e-8 k1=0.64774 k2=6.160789912e-02 wk2=-2.046758304e-8 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=123760.0 ua=-3.385286549e-09 wua=1.824486888e-16 ub=3.462877957e-18 wub=-2.008450572e-25 uc=1.321115660e-11 wuc=2.484375444e-17 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=9.678542589e-04 wu0=6.013015329e-10 a0=2.543343285e+00 wa0=-5.118518969e-7 keta=-0.01258 a1=0.0 a2=0.46703705 ags=7.229106026e-01 wags=-2.420312796e-7 b0=5.217906632e-07 wb0=-1.945470064e-13 b1=4.764694966e-07 wb1=-1.444006705e-13 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-5.732703382e-02+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' wvoff=-5.455778509e-8 nfactor='2.065275749e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' wnfactor=2.603151055e-7 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-5.291112804e-01 wpclm=3.351883249e-7 pdiblc1=0.0 pdiblc2=5.465828918e-03 wpdiblc2=1.016561674e-9 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.914848965e-02 wdelta=-2.755126701e-9 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-6.685948551e-01 wkt1=-8.999070560e-8 kt2=-0.055045 at=232120.0 ute=-4.041480806e-02 wute=-3.316540579e-8 ua1=6.9609e-10 ub1=-1.2188e-19 uc1=-9.961e-12 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=3.0e-6 sbref=3.0e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.45 pmos lmin=1e-06 lmax=1.5e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='1.426706620e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=-3.385230616e-07 wvth0=-2.018771487e-07 pvth0=1.989632040e-13 k1=0.64774 k2=1.294794950e-01 lk2=-9.907556202e-08 wk2=-7.346856138e-08 pk2=7.736817814e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=3.918191587e+05 lvsat=-3.912993570e-01 wvsat=-1.258264330e-01 pvsat=1.836751356e-7 ua=-4.576715022e-09 lua=1.739187714e-15 wua=5.368132799e-16 pua=-5.172837118e-22 ub=5.345945005e-18 lub=-2.748807124e-24 wub=-9.423934688e-25 pub=1.082475294e-30 uc=-8.966149132e-11 luc=1.501683478e-16 wuc=6.535265394e-17 puc=-5.913286605e-23 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=-3.530444769e-04 lu0=1.928181930e-09 wu0=6.391973570e-10 pu0=-5.531842930e-17 a0=4.686504709e+00 la0=-3.128479890e-06 wa0=-1.369721628e-06 pa0=1.252275340e-12 keta=-7.470874428e-02 lketa=9.069243446e-08 wketa=3.637118399e-08 pketa=-5.309283584e-14 a1=0.0 a2=0.46703705 ags=-9.927243005e-01 lags=2.504398050e-06 wags=6.127227017e-07 pags=-1.247727124e-12 b0=-3.919334347e-07 lb0=1.333808752e-12 wb0=1.932059577e-13 pb0=-5.660223893e-19 b1=5.193923699e-07 lb1=-6.265666425e-14 wb1=-3.079982976e-13 pb1=2.388116362e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='1.485152689e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-3.004783014e-07 wvoff=-1.994164631e-07 pvoff=2.114574552e-13 nfactor='3.464220939e-01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.509096623e-06 wnfactor=1.273561039e-06 pnfactor=-1.479085751e-12 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-5.291112804e-01 wpclm=3.351883249e-7 pdiblc1=0.0 pdiblc2=-4.715720763e-02 lpdiblc2=7.681647760e-08 wpdiblc2=1.757033173e-08 ppdiblc2=-2.416436584e-14 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=2.099183397e-02 ldelta=1.190667812e-08 wdelta=-5.704703016e-09 pdelta=4.305644026e-15 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-1.013593083e-01 lkt1=-8.280220895e-07 wkt1=-4.269070987e-07 pkt1=4.918137049e-13 kt2=3.104333000e-03 lkt2=-8.488348885e-8 at=1.027896501e+06 lat=-1.161634747e+00 wat=-3.372071964e-01 pat=4.922382050e-7 ute=-1.894130284e-01 lute=2.175001522e-07 wute=6.103824564e-08 pute=-1.375137802e-13 ua1=3.433807053e-10 lua1=5.148673930e-16 wua1=1.802565018e-16 pua1=-2.631294285e-22 ub1=-4.880210018e-19 lub1=5.344743274e-25 wub1=1.873271763e-25 pub1=-2.734508456e-31 uc1=-8.666613950e-11 luc1=1.119703274e-16 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=2.74e-6 sbref=2.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.46 pmos lmin=5e-07 lmax=1e-06 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-1.721325756e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))' lvth0=-3.639065436e-08 wvth0=-2.646044352e-08 pvth0=3.060702122e-14 k1=0.64774 k2=3.724395733e-02 lk2=-1.055250478e-08 wk2=5.174130109e-09 pk2=1.890854977e-15 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=1.523299471e+05 lvsat=-1.614495861e-01 wvsat=-2.123061246e-02 pvsat=8.328929680e-8 ua=-2.778837784e-09 lua=1.367503439e-17 wua=8.221401961e-17 pua=-8.098207174e-23 ub=2.092687198e-18 lub=3.735070566e-25 wub=2.599067061e-25 pub=-7.143229913e-32 uc=8.813146605e-11 luc=-2.046844304e-17 wuc=-6.061143475e-18 puc=9.406526022e-24 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=1.081899490e-03 lu0=5.509944573e-10 wu0=1.018013691e-09 pu0=-4.188874059e-16 a0=3.418373795e+00 la0=-1.911391245e-06 wa0=-1.172791534e-06 pa0=1.063271682e-12 keta=4.634785522e-02 lketa=-2.549163690e-08 wketa=-3.486869307e-08 pketa=1.527963618e-14 a1=0.0 a2=0.46703705 ags=1.489515562e+00 lags=1.220683421e-07 wags=-6.276299824e-07 pags=-5.729863566e-14 b0=1.392972995e-06 lb0=-3.792551938e-13 wb0=-5.796730989e-13 pb0=1.757482853e-19 b1=-5.551016968e-08 lb1=4.891060481e-13 wb1=2.309984256e-13 pb1=-2.784904689e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='-1.697816508e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=5.007167319e-09 wvoff=2.451905421e-08 pvoff=-3.464657503e-15 nfactor='2.728110446e+00+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=2.232712266e-07 wnfactor=-5.526160525e-08 pnfactor=-2.037482186e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=0.0 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-9.344276432e-01 lpclm=3.890023792e-07 wpclm=5.781341421e-07 ppclm=-2.331672481e-13 pdiblc1=0.0 pdiblc2=-1.273572964e-01 lpdiblc2=1.537885128e-07 wpdiblc2=5.707927250e-08 ppdiblc2=-6.208307174e-14 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=9.972205229e-02 ldelta=-6.365464891e-08 wdelta=-4.269320853e-08 pdelta=3.980536220e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-2.668682491e-01 lkt1=-6.691748835e-07 wkt1=-7.367204470e-08 pkt1=1.527963618e-13 kt2=-0.085339 at=-3.552405265e+05 lat=1.658310149e-01 wat=2.849682736e-01 pat=-1.048947024e-7 ute=1.633719963e-01 lute=-1.210852753e-07 wute=-1.578646478e-07 pute=7.257827184e-14 ua1=9.278490842e-10 lua1=-4.607613370e-17 wua1=-1.226842337e-16 pua1=2.761794239e-23 ub1=9.513846034e-19 lub1=-8.469952022e-25 wub1=-5.246015628e-25 pub1=4.098227617e-31 uc1=3.0e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.74e-6 sbref=1.74e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.model sky130_fd_pr__pfet_01v8_lvt__model.47 pmos lmin=3.5e-07 lmax=5e-07 wmin=4.2e-07 wmax=5.5e-7 level=54.0 tnom=30.0 version=4.5 toxm=4.23e-9 xj=1.5e-7 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint=2.0125e-8 ll=0.0 lw=0.0 lwl=0.0 wint=-2.4699e-8 wl=0.0 ww=0.0 wwl=0.0 xl=0.0 xw=0.0 mobmod=0.0 binunit=2.0 dwg=-7.916e-9 dwb=0.0 igcmod=0.0 igbmod=0.0 rgatemod=0.0 rbodymod=1.0 trnqsmod=0.0 acnqsmod=0.0 fnoimod=1.0 tnoimod=1.0 permod=1.0 geomod=0.0 rdsmod=0.0 tempmod=0.0 lintnoi=0.0 vfbsdoff=0.0 lambda=0.0 vtl=0.0 lc=5.0e-9 xn=3.0 rnoia=0.69 rnoib=0.34 tnoia=25000000.0 tnoib=0.0 epsrox=3.9 toxe='4.01004e-09+sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre*(4.01004e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))' dtox=0.0 ndep=1.7000000000000000e+17 nsd=1.0e+20 rshg=0.1 rsh=1.0 vth0='-3.591445216e-01+sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))' lvth0=4.958808782e-08 wvth0=-1.662867217e-08 pvth0=2.608686434e-14 k1=0.64774 k2=-5.783588913e-02 lk2=3.316045463e-08 wk2=-1.864133227e-08 pk2=1.284001380e-14 k3=3.39 dvt0=2.4422 dvt1=0.16136 dvt2=0.026237 dvt0w=0.5 dvt1w=1928100.0 dvt2w=-0.032 w0=1.0e-8 k3b=1.0 phin=0.0 lpe0=0.0 lpeb=0.0 vbm=-3.0 dvtp0=0.0 dvtp1=0.0 vsat=-4.317216670e+05 lvsat=1.070681435e-01 wvsat=2.375085216e-01 pvsat=-3.566602010e-8 ua=-2.061790088e-09 lua=-3.159876438e-16 wua=-3.576145801e-16 pua=1.212291270e-22 ub=1.317011342e-18 lub=7.301240316e-25 wub=7.239706815e-25 pub=-2.847857118e-31 uc=7.453845146e-11 luc=-1.421905458e-17 wuc=8.521901228e-18 puc=2.701971220e-24 rdsw=484.7 prwb=0.1 prwg=0.052 wr=1.0 u0=3.582810484e-03 lu0=-5.987993722e-10 wu0=-2.039010187e-11 pu0=5.851873790e-17 a0=-7.390840508e-01 wa0=1.139925556e-6 keta=-9.098880846e-03 wketa=-1.634030369e-9 a1=0.0 a2=0.46703705 ags=4.240346405e+00 lags=-1.142626138e-06 wags=-1.918864479e-06 pags=5.363464239e-13 b0=1.741094271e-06 lb0=-5.393039504e-13 wb0=-6.050428131e-13 pb0=1.874120114e-19 b1=3.090568317e-06 lb1=-9.573035363e-13 wb1=-1.148592951e-12 pb1=3.557766667e-19 eu=1.67 rdswmin=0.0 rdw=0.0 rdwmin=0.0 rsw=0.0 rswmin=0.0 voff='8.178738557e-01+sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))' lvoff=-4.490674518e-07 wvoff=5.205318446e-08 pvoff=-1.612347389e-14 nfactor='-1.190939114e+01+sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))' lnfactor=6.952862580e-06 wnfactor=-1.527698277e-06 pnfactor=4.732045413e-13 up=0.0 ud=0.0 lp=1.0 tvfbsdoff=0.0 tvoff=4.473724015e-2 cit=-6.393105e-11 cdsc=2.8125e-7 cdscb=1.0e-4 cdscd=1.0e-10 eta0=0.2 etab=-0.00025 dsub=1.0 voffl=0.0 minv=0.0 pclm=-8.831045088e-02 wpclm=7.097318924e-8 pdiblc1=0.0 pdiblc2=-4.564133840e-02 lpdiblc2=1.162196011e-07 wpdiblc2=-1.469082037e-08 ppdiblc2=-2.908677155e-14 pdiblcb=-0.025 drout=4.663735585e-01 wdrout=-1.882922411e-8 pscbe1=800000000.0 pscbe2=8.6797e-9 pvag=0.0 delta=1.249506561e-01 ldelta=-7.525349952e-08 wdelta=-5.736328537e-08 pdelta=4.654993002e-14 alpha0=5.0449517e-13 alpha1=-4.0583656e-18 beta0=6.2016506 fprout=0.0 pdits=0.0 pditsl=0.0 pditsd=0.0 agidl=0.0 bgidl=2300000000.0 cgidl=0.5 egidl=0.8 aigbacc=0.43 bigbacc=0.054 cigbacc=0.075 nigbacc=1.0 aigbinv=0.35 bigbinv=0.03 cigbinv=0.006 eigbinv=1.1 nigbinv=3.0 aigc=0.43 bigc=0.054 cigc=0.075 nigc=1.0 aigsd=0.43 bigsd=0.054 cigsd=0.075 dlcig=0.0 poxedge=1.0 pigcd=1.0 ntox=1.0 toxref=4.23e-9 kt1=-5.916684453e+00 lkt1=1.928328116e-06 wkt1=2.795725430e-06 pkt1=-1.166409127e-12 kt2=-0.085339 at=-5.123944135e+03 lat=4.864916196e-03 wat=1.741297428e-01 pat=-5.393668784e-8 ute=1.320027500e-01 lute=-1.066632643e-07 pute=2.524354897e-29 ua1=1.043337168e-09 lua1=-9.917178040e-17 wua1=-1.919075604e-16 pua1=5.944336683e-23 ub1=-2.250590322e-18 lub1=6.251127698e-25 wub1=1.124247955e-24 pub1=-3.482358040e-31 uc1=3.0e-11 kt1l=0.0 prt=0.0 xrcrg1=12.0 xrcrg2=1.0 rbpb=50.0 rbpd=50.0 rbps=50.0 rbdb=50.0 rbsb=50.0 gbmin=1.0e-12 noia=3.0e+41 noib=0.0 noic=0.0 em=41000000.0 af=1.0 ef=0.88 kf=0.0 ntnoi=1.0 dmcg=0.0 dmcgt=0.0 dmdg=0.0 xgw=0.0 xgl=0.0 ngcon=1.0 diomod=1.0 njs=1.3632 jss=2.1483e-5 jsws=1.4472e-10 xtis=5.2 bvs=12.69 xjbvs=1.0 ijthsrev=0.1 ijthsfwd=0.1 tpb=0.001671 tpbsw=0.001246 tpbswg=0.0 tcj=0.0012407 tcjsw=0.00037357 tcjswg=2.0e-12 cgdo=1.0e-11 cgso=1.0e-11 cgbo=1.0e-13 capmod=2.0 xpart=0.0 cgsl=0.0 cgdl=0.0 cf=0.0 clc=7.0e-8 cle=0.492 dlc=3.417e-8 dwc=-3.2175e-8 vfbcv=-1.0 acde=0.44 moin=8.7 noff=2.6123 voffcv=0.112 ngate=1.0e+23 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 ckappas=0.6 cjs=0.0006926438503 mjs=0.3362 pbs=0.6587 cjsws=8.29052224e-11 mjsws=0.2659 pbsws=0.7418 cjswgs=2.164485778e-10 mjswgs=0.9274 pbswgs=1.4338 saref=1.44e-6 sbref=1.44e-6 wlod='0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff' kvth0='0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff' lkvth0='0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff' wkvth0='0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff' pkvth0=0.0 llodvth=0.0 wlodvth=1.0 stk2=0.0 lodk2=1.0 lodeta0=1.0 ku0='0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff' lku0='0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff' wku0='0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff' pku0=0.0 llodku0=0.0 wlodku0=1.0 kvsat='0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff' steta0=0.0 tku0=0.0
.ends sky130_fd_pr__pfet_01v8_lvt