* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.subckt sky130_fd_pr__res_xhigh_po_0p35 r0 r1 b
.param w=0.35
.param l=5
.param mult=1.0
xsky130_fd_pr__res_xhigh_po_0p35 r0 r1 b sky130_fd_pr__res_xhigh_po__base w='w' l='l' mult='mult'
.ends sky130_fd_pr__res_xhigh_po_0p35