* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__res_high_po__var_mult=5.0
.param sky130_fd_pr__res_high_po__var=0.125
.param sky130_fd_pr__res_xhigh_po__var_mult=0.15
.param camimc=1.778e-15
.param cpmimc=0.03e-15
.param cvpp_cor=0.862
.param cvpp3_cor=0.7
.param cvpp4_cor=0.7
.param cvpp5_cor=0.7
.param cm3m2_vpp=0.446
.param c0m5m4_vpp=0.804
.param c1m5m4_vpp=0.766
.param c0m5m4_vpp0p4shield=0.6046
.param c1m5m4_vpp0p4shield=0.766
.param c0m4m3_vpp=0.804
.param c1m4m3_vpp=0.766
.param c0m5m3_vpp=0.803
.param c1m5m3_vpp=0.774
.param cpl2s_vpp=0.760
.param cpl2s_vpp0p4shield=0.7511
.param cli2s_vpp=0.794
.param sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1__cor=0.810
.param sky130_fd_pr__cap_vpp_04p4x04p6_m1m2m3_shieldl1__cor=0.775
.param sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3_shieldl1__cor=0.855
.param sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield__cor=0.827
.param sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield__cor=0.796
.param sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield__cor=0.868
.param sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield__cor=0.786
.param sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1__cor=0.827
.param sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1__cor=0.796
.param sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1__cor=0.868
.param sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3__cor=0.846
.param sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3__cor=0.816
.param sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3__cor=0.885
.param sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3__cor=0.863
.param sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5__cor=0.856
.param sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldpom5__cor=0.856
.param sky130_fd_pr__cap_vpp_11p5x11p7_m1m2m3m4_shieldl1m5__cor=0.856
.param sky130_fd_pr__cap_vpp_08p6x07p8_m1m2m3_shieldl1m5_floatm4__cor=0.792
.param sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2_noshield__cor=0.8
.param sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldm4__cor=0.8
.param sky130_fd_pr__model__cap_vpp_finger__cor=0.8
.param sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield_base__cor=0.8