* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_pfet_01v8_b__toxe_mult=0.9635
.param sky130_fd_pr__rf_pfet_01v8_b__rbpb_mult=0.8
.param sky130_fd_pr__rf_pfet_01v8_b__overlap_mult=0.88516
.param sky130_fd_pr__rf_pfet_01v8_b__ajunction_mult=0.93001
.param sky130_fd_pr__rf_pfet_01v8_b__pjunction_mult=0.93439
.param sky130_fd_pr__rf_pfet_01v8_b__lint_diff=1.21275e-8
.param sky130_fd_pr__rf_pfet_01v8_b__wint_diff=-2.252e-8
.param sky130_fd_pr__rf_pfet_01v8_b__rshg_diff=-7.0
.param sky130_fd_pr__rf_pfet_01v8_b__dlc_diff=1.21275e-8
.param sky130_fd_pr__rf_pfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_pfet_01v8_b__xgw_diff=-4.504e-8
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult=0.8875
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult=0.839
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult=0.839
.param sky130_fd_pr__rf_pfet_01v8__aw_cap_mult_2=0.8875
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_dist_mult_2=0.86
.param sky130_fd_pr__rf_pfet_01v8__aw_rgate_stub_mult_2=0.86
.param sky130_fd_pr__rf_pfet_01v8__aw_rd_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8__aw_rs_mult=1.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_0=-0.0096187
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_0=-9.1722e-5
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_0=-0.057483
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_0=-11003.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_1=-0.012861
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_1=1.6284e-5
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_1=-0.054689
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_1=-6396.5
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_2=-0.029824
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_2=0.00016037
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_2=-0.02191
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_2=5271.4
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_3=-0.013607
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_3=3.7455e-6
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_3=-0.077102
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_3=-10440.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_4=-0.0077158
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_4=-0.00015599
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_4=-0.04551
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_4=-2665.7
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_5=-0.018523
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_5=2.6323e-5
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_5=-0.017911
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_5=11962.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_6=-0.013977
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_6=-0.00029174
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_6=-0.081869
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_6=-8538.5
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_7=-3.0985e-5
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_7=-8661.9
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_7=-0.0068507
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_7=-0.050877
.param sky130_fd_pr__rf_pfet_01v8_bm02__vth0_diff_8=-0.024781
.param sky130_fd_pr__rf_pfet_01v8_bm02__u0_diff_8=-3.1187e-5
.param sky130_fd_pr__rf_pfet_01v8_bm02__vsat_diff_8=3310.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm02__k2_diff_8=-0.020378
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_0=-0.007218
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_0=-0.00024908
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_0=-0.045584
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_0=-10840.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_1=-0.011746
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_1=-5.8756e-5
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_1=-0.040864
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_1=-2721.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_2=0.00011377
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_2=-0.014596
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_2=11806.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_2=-0.030918
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_3=-0.011489
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_3=-0.00010472
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_3=-0.075251
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_3=-6951.2
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_4=-0.00033553
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_4=-0.032126
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_4=-3166.2
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_4=-0.0039733
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_5=-0.0099782
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_5=-7.0926e-5
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_5=7638.8
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_5=-0.018384
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_6=-0.076598
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_6=-0.00010558
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_6=-8165.2
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_6=-0.012381
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_7=-0.0043219
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_7=-0.046792
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_7=-0.00030508
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_7=-6293.3
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__k2_diff_8=-0.018996
.param sky130_fd_pr__rf_pfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vth0_diff_8=-0.012116
.param sky130_fd_pr__rf_pfet_01v8_bm04__u0_diff_8=-0.00013862
.param sky130_fd_pr__rf_pfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__vsat_diff_8=17138.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_pfet_01v8_bm04__ub_diff_8=0.0
.include "sky130_fd_pr__rf_pfet_01v8_b.pm3.spice"