* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param tol_nfom=0.0483u
.param tol_pfom=0.042u
.param tol_nw=0.0483u
.param tol_poly=0.0287u
.param tol_li=0.014u
.param tol_m1=0.0175u
.param tol_m2=0.0175u
.param tol_m3=0.0455u
.param tol_m4=0.0455u
.param tol_m5=0.119u
.param tol_rdl=0.7u
.param rcn=103.6
.param rcp=411
.param rdn=111.6
.param rdp=175.3
.param rdn_hv=105.6
.param rdp_hv=169.3
.param rp1=44
.param rnw=1378
.param rl1=10.31
.param rm1=0.111
.param rm2=0.111
.param rm3=0.0407
.param rm4=0.0407
.param rm5=0.02339
.param rrdl=0.0043
.param rcp1=61.28
.param rcl1=3.91
.param rcvia=2.75
.param rcvia2=1.373
.param rcvia3=1.373
.param rcvia4=0.1224
.param rcrdlcon=0.00496
.param rspwres=3512
.param crpf_precision=8.84e-5
.param crpfsw_precision_1_1=4.67e-11
.param crpfsw_precision_2_1=5.02e-11
.param crpfsw_precision_4_1=5.45e-11
.param crpfsw_precision_8_2=5.96e-11
.param crpfsw_precision_16_2=6.54e-11
.include "../sky130_fd_pr__model__r+c.model.spice"
.include "../parameters/fast_70p.spice"