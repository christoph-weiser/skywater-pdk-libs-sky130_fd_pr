* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__special_nfet_latch__tox_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_latch__vth0_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_latch__voff_slope_spectre=0.0
.param sky130_fd_pr__special_nfet_latch__nfactor_slope_spectre=0.0
.subckt sky130_fd_pr__special_nfet_latch d g s b
.param l=1
.param w=1
.param ad=0
.param as=0
.param pd=0
.param ps=0
.param nrd=0
.param nrs=0
.param mult=1
.param sa=0
.param sb=0
.param sd=0.0
msky130_fd_pr__special_nfet_latch d g s b sky130_fd_pr__special_nfet_latch__model l='l' w='w' ad='ad' as='as' pd='pd' ps='ps' nrd='nrd' nrs='nrs'
.model sky130_fd_pr__special_nfet_latch__model.0 nmos lmin=7.5e-08 lmax=1.505e-007 wmin=2.095e-007 wmax=2.105e-7 level=49.0 tnom=30.0 version=3.2 tox='4.148e-009*sky130_fd_pr__special_nfet_latch__tox_mult+sky130_fd_pr__special_nfet_latch__tox_slope_spectre*(4.148e-009*sky130_fd_pr__special_nfet_latch__tox_mult*(sky130_fd_pr__special_nfet_latch__tox_slope/sqrt(l*w*mult)))' toxm=4.148e-9 xj=1.2e-7 nch=1.12471e+18 lln=1.0 lwn=1.0 wln=1.0 wwn=1.0 lint='0+sky130_fd_pr__special_nfet_latch__lint_diff' ll=0.0 lw=0.0 lwl=0.0 wint='0+sky130_fd_pr__special_nfet_latch__wint_diff' wl=0.0 ww=0.0 wwl=0.0 mobmod=1.0 binunit=2.0 dwg=0.0 dwb=0.0 ldif=0.0 hdif=0.0 rd=0.0 rs=0.0 rsc=0.0 rdc=0.0 rsh=1.0 vth0='0.71908+sky130_fd_pr__special_nfet_latch__vth0_diff_0+sky130_fd_pr__special_nfet_latch__vth0_slope_spectre*(sky130_fd_pr__special_nfet_latch__vth0_slope/sqrt(l*w*mult))' k1=0.498 k2='-0.1068+sky130_fd_pr__special_nfet_latch__k2_diff_0' k3='0+sky130_fd_pr__special_nfet_latch__k3_diff' dvt0='0+sky130_fd_pr__special_nfet_latch__dvt0_diff' dvt1='0.53+sky130_fd_pr__special_nfet_latch__dvt1_diff' dvt2=0.0 dvt0w=0.0 dvt1w=0.0 dvt2w=0.0 nlx=0.0 w0=0.0 k3b=0.0 ngate=1.0e+23 vfb=-0.9693 vsat='82072+sky130_fd_pr__special_nfet_latch__vsat_diff_0' ua=-1.048e-9 ub=1.2106e-18 uc=6.2252e-11 rdsw='187.1195+sky130_fd_pr__special_nfet_latch__rdsw_diff_0' prwb=0.3 prwg=0.2 wr=1.0 u0='0.022616+sky130_fd_pr__special_nfet_latch__u0_diff_0' a0=-0.1 keta=-0.019632 a1=0.0 a2=0.99 ags=0.02 b0=0.0 b1=0.0 voff='-0.139+sky130_fd_pr__special_nfet_latch__voff_diff_0+sky130_fd_pr__special_nfet_latch__voff_slope_spectre*(sky130_fd_pr__special_nfet_latch__voff_slope/sqrt(l*w*mult))' nfactor='1.078+sky130_fd_pr__special_nfet_latch__nfactor_diff_0+sky130_fd_pr__special_nfet_latch__nfactor_slope_spectre*(sky130_fd_pr__special_nfet_latch__nfactor_slope/sqrt(l*w*mult))' cit='0+sky130_fd_pr__special_nfet_latch__cit_diff' cdsc='0+sky130_fd_pr__special_nfet_latch__cdsc_diff' cdscb='0+sky130_fd_pr__special_nfet_latch__cdscb_diff' cdscd='0+sky130_fd_pr__special_nfet_latch__cdscd_diff' eta0=0.01 etab=-0.0042 dsub=0.0 pclm=0.9345125 pdiblc1=0.0 pdiblc2=0.024526 pdiblcb=0.05573667 drout=0.0 pscbe1=7.7384e+8 pscbe2=9.2e-21 pvag=0.0 delta=0.023 alpha0=4.1e-6 alpha1=0.0 beta0=17.69 kt1='-0.2357+sky130_fd_pr__special_nfet_latch__kt1_diff_0' kt2='-0.02+sky130_fd_pr__special_nfet_latch__kt2_diff' at=31512.0 ute=-1.25 ua1=5.5e-10 ub1=-2.0e-19 uc1=-3.5e-12 kt1l=0.0 prt=-8.0505 cj='0.0013459*sky130_fd_pr__special_nfet_latch__ajunction_mult' mj=0.44 pb=0.729 cjsw='3.6001e-011*sky130_fd_pr__special_nfet_latch__pjunction_mult' mjsw=0.0009 pbsw=0.2 cjswg='2.3347e-010*sky130_fd_pr__special_nfet_latch__pjunction_mult' mjswg=0.8000 pbswg=0.95578 tpb=0.0012287 tpbsw=0.0 tpbswg=0.0 tcj=0.000792 tcjsw=1.0e-5 tcjswg=0.0 js=0.0027500000000000003 jsw=6.0e-10 nj=1.2928 xti=2.0 cgdo='3.2e-010*sky130_fd_pr__special_nfet_latch__overlap_mult' cgso='3.2e-010*sky130_fd_pr__special_nfet_latch__overlap_mult' cgbo=1.0e-13 capmod=3.0 nqsmod=0.0 elm=0.0 xpart=0.0 cgsl='0*sky130_fd_pr__special_nfet_latch__overlap_mult' cgdl='0*sky130_fd_pr__special_nfet_latch__overlap_mult' ckappa=0.6 cf=1.4067e-12 clc=1.0e-7 cle=0.6 dlc='1.8739e-008+sky130_fd_pr__special_nfet_latch__dlc_diff+sky130_fd_pr__special_nfet_latch__dlc_rotweak' dwc='0+sky130_fd_pr__special_nfet_latch__dwc_diff' vfbcv=-1.0 acde=0.4 moin=6.9 noff=3.621 voffcv=-0.1372 lwc=0.0 llc=0.0 lwlc=0.0 wlc=0.0 wwc=0.0 wwlc=0.0 noimod=2.0 noia='1.1737146e+41*1.6e-21' noib='3.2036721e+25*1.6e-21' noic='-3.7339643e+08*1.6e-21' em=4.1000000e+7 ef=0.8439365
.ends sky130_fd_pr__special_nfet_latch