* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.model sky130_fd_pr__diode_pw2nd_05v5_nvt d level=3.0 tlevc=1.0 area=1.0e+12 cj='0.0008602*1e-12*sky130_fd_pr__nfet_05v0_nvt__ajunction_mult' mj=0.28329 pb=0.66345 cjsw='8.5152e-011*1e-6*sky130_fd_pr__nfet_05v0_nvt__pjunction_mult' mjsw=0.057926 php=1 cta=0.00083 ctp=0 tpb=0.0019685 tphp=0.001 js=4.2966e-016 jsw=8.04e-016 n=1.5764 rs=600 ik='4.76e-008/1e-12' ikr='0/1e-12' vb=12.69 ibv=0.00106 trs=0 eg=1.05 xti=0.0 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0