* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param ndiodedefet_pb_mult=2.7281
.model sky130_fd_pr__diode_pw2nd_05v5__extended_drain d level=3.0 tlevc=1.0 scalm=1.0e-6 area=1.0e+12 cj='0.0013459*1e-12*sky130_fd_pr__nfet_01v8__ajunction_mult' mj=0.44 pb='0.729*ndiodedefet_pb_mult' cjsw='3.6001e-011*1e-6*sky130_fd_pr__nfet_01v8__pjunction_mult' mjsw=0.0009 php=0.2 cta=0.000792 ctp=1e-005 tpb=0.0012287 tphp=0 js=2.75e-015 jsw=6e-016 n=1.2928 rs=981 ik='1.3e-009/1e-12' ikr='0/1e-12' vb=11.7 ibv=0.00106 trs=0 eg=1.05 xti=2.0 tref=30 tcv=0 gap1=0.000473 gap2=1110.0 ttt1=0 ttt2=0 tm1=0 tm2=0 lm=0 lp=0 wm=0 wp=0 xm=0 xoi=10000.0 xom=10000 xp=0 xw=0