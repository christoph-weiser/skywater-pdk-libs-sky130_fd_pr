* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param dkisnpn1x1=8.7913e-01
.param dkbfnpn1x1=9.8501e-01
.param dkisnpn1x2=9.0950e-01
.param dkbfnpn1x2=9.6759e-01
.param dkisnpnpolyhv=1.0
.param dkbfnpnpolyhv=1.0
.include "sky130_fd_pr__npn_05v5_W1p00L1p00.model.spice"
.include "sky130_fd_pr__npn_05v5_W1p00L2p00.model.spice"
.include "../npn_11v0/sky130_fd_pr__npn_11v0_W1p00L1p00.model.spice"