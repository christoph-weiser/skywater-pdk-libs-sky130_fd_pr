* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_20v0__toxe_mult=0.94
.param sky130_fd_pr__nfet_20v0__rshn_mult=1.0
.param sky130_fd_pr__nfet_20v0__overlap_mult=1.9
.param sky130_fd_pr__nfet_20v0__ajunction_mult=4.1753e-1
.param sky130_fd_pr__nfet_20v0__pjunction_mult=4.7786e-1
.param sky130_fd_pr__nfet_20v0__lint_diff=1.7325e-8
.param sky130_fd_pr__nfet_20v0__wint_diff=-3.2175e-8
.param sky130_fd_pr__nfet_20v0__dlc_diff=1.7325e-8
.param sky130_fd_pr__nfet_20v0__dwc_diff=-3.2175e-8
.param sky130_fd_pr__nfet_20v0__rdrift_mult=4.9875e-1
.param sky130_fd_pr__nfet_20v0__hvvsat_mult=5.6124e-1
.param sky130_fd_pr__nfet_20v0__vth0_diff=-1.0850e-1
.param sky130_fd_pr__nfet_20v0__k2_diff=-2.8999e-2
.param sky130_fd_pr__nfet_20v0_iso__rdrift_mult=2.8388e-1
.param sky130_fd_pr__nfet_20v0_iso__hvvsat_mult=2.1534e-1
.param sky130_fd_pr__nfet_20v0_iso__vth0_diff=-1.4327e-1
.param sky130_fd_pr__nfet_20v0_iso__k2_diff=-2.0083e-2
.include "sky130_fd_pr__nfet_20v0__subcircuit.pm3.spice"
.include "../nfet_20v0_iso/sky130_fd_pr__nfet_20v0_iso__subcircuit.pm3.spice"
.include "../nfet_20v0_zvt/sky130_fd_pr__nfet_20v0_zvt__sf_discrete.corner.spice"