* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_lvt__toxe_slope=6.789e-03
.param sky130_fd_pr__rf_nfet_01v8_lvt__toxe1_slope=8.089e-03
.param sky130_fd_pr__rf_nfet_01v8_lvt__b_toxe_slope=3.443e-03
.param sky130_fd_pr__rf_nfet_01v8_lvt__b_vth0_slope=6.056e-03