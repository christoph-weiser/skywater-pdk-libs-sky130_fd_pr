* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__pfet_g5v0d10v5__toxe_mult=0.94
.param sky130_fd_pr__pfet_g5v0d10v5__rshp_mult=1.0
.param sky130_fd_pr__pfet_g5v0d10v5__overlap_mult=0.7
.param sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult=0.93222
.param sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult=0.94436
.param sky130_fd_pr__pfet_g5v0d10v5__lint_diff=1.7325e-8
.param sky130_fd_pr__pfet_g5v0d10v5__wint_diff=-3.2175e-8
.param sky130_fd_pr__pfet_g5v0d10v5__dlc_diff=1.7325e-8
.param sky130_fd_pr__pfet_g5v0d10v5__dwc_diff=-3.2175e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0=7.1446e-9
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0=-8.1068e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0=-5.8946e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0=0.0023082
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0=0.019265
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0=0.78564
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0=-0.0024588
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0=0.026115
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0=-3965.1
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1=6.7197e-9
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1=-1.0086e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1=1.3345e-12
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1=0.074623
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1=-0.021649
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1=0.0080331
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1=2.4188
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1=-0.00091756
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1=0.10857
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1=-0.034924
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2=1.1489e-8
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2=-6.4117e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2=2.5554e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2=0.023145
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2=0.020797
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2=0.64494
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2=-0.0021939
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2=0.046498
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2=-3087.7
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3=-0.069521
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3=7.4686e-9
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3=-3.3536e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3=2.7072e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3=-0.20155
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3=0.026441
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3=0.0032184
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3=2.0168
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3=-0.0012151
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3=0.095591
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4=2.4859
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4=-0.00096391
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4=0.098544
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4=-0.031072
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4=1.023e-8
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4=-3.0365e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4=-1.9852e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4=-0.28336
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4=0.0069066
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4=0.0026716
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5=-0.1047086
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5=3.5856
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5=-0.0018767
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5=0.14168
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5=0.0028699
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5=0.00016238
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5=2.3237e-8
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5=-5.045e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5=1.2416e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5=-0.12955
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5=-0.0002908
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6=0.019041
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6=0.84301
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6=-0.0034483
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6=0.076423
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6=-9946.4
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6=3.9908e-8
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6=-1.1687e-18
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6=-2.1854e-12
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6=0.030875
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7=-0.023831
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7=0.0084689
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7=0.092518
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7=1.67
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7=-0.0013725
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7=-0.047184
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7=-1.5753e-10
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7=-4.2337e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7=-3.5098e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7=-0.12601
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8=-0.19863
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8=-0.032394
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8=0.0067604
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8=0.12076
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8=2.4084
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8=-0.0014593
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8=-0.053538
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8=1.4663e-7
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8=-5.0813e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8=-5.8602e-13
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9=-0.38314
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9=0.0047331
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9=0.0025401
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9=0.1075
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9=2.8659
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9=-0.0010746
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9=-0.025322
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9=1.6873e-7
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9=-2.6015e-19
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9=-2.9672e-14
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10=1.49e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10=3.7525
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10=-0.0010652
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10=-0.26081
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10=0.14547
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10=-0.015852
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10=0.0033082
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10=3.7574e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10=-1.9776e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10=0.0074642
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10=0.0022763
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11=-20938.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11=9.5411e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11=0.39133
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11=-0.0019065
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11=0.076426
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11=0.022745
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11=0.019312
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11=8.5779e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11=-4.1882e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12=-9517.3
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12=1.1957e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12=1.3162
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12=-0.0031096
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12=0.022012
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12=0.097785
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12=0.011937
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12=-8.4463e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12=-8.4748e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13=-6.9753e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13=0.0012324
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13=-4426.9
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13=2.2526e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13=1.4877
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13=-0.002059
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13=-0.065209
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13=0.083581
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13=0.012626
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13=-1.3471e-12
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14=6.5821e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14=-4.0194e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14=-0.016665
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14=8.3957e-10
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14=2.4556
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14=-0.0015647
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14=0.068222
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14=0.1083
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14=-0.026998
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14=0.008511
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15=0.018378
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15=3.9683e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15=-7.8901e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15=-3884.3
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15=-1.4078e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15=0.93444
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15=-0.0027952
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15=0.018219
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15=0.028672
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16=-0.064881
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16=0.098497
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16=-0.030763
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16=0.008808
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16=4.6538e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16=-6.6411e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16=0.0011356
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16=-0.016503
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16=8.1848e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16=1.991
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16=-0.0025485
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17=1.365e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17=3.2265
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17=-0.00068848
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17=-0.00048569
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17=0.11349
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17=-0.013211
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17=0.0016068
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17=1.4383e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17=1.57e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17=0.0015256
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18=1.3923e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18=3.305
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18=-0.0021335
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18=-0.37258
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18=0.12843
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18=-0.0095856
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18=0.0029978
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18=4.4933e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18=-5.6175e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18=0.0018439
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19=5.8126e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19=3.2747
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19=-0.0014519
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19=-0.17225
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19=0.13332
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19=-0.0050121
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19=0.00066506
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19=6.1444e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19=-3.157e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19=0.0059198
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19=0.00066294
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20=1.0061e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20=1.0343
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20=-0.0021126
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20=0.021271
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20=0.027094
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20=0.020516
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20=1.4571e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20=-4.573e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20=-23962.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21=-7800.3
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21=2.3024e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21=1.0441
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21=-0.0032065
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21=0.16212
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21=0.076409
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21=0.015471
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21=-5.568e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21=-8.928e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22=-0.010622
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22=-0.030587
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22=-2.6823e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22=1.9965
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22=-0.00011051
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22=-0.13262
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22=0.057087
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22=-0.017178
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22=0.0040145
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22=2.3221e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22=2.4278e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23=0.00021003
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23=5.5063e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23=2.5904
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23=-0.0011579
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23=-0.24208
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23=0.084349
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23=-0.0037978
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23=0.00031172
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23=1.2987e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23=-2.3608e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24=-6.3305e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24=0.0010943
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24=2.7509e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24=3.4168
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24=-0.0025093
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24=-0.29695
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24=0.12799
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24=-0.0034495
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24=0.0035991
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24=8.8967e-13
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25=8.0711e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25=-5.0441e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25=-0.00085579
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25=-1.069e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25=3.4716
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25=-0.002061
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25=-0.26818
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25=0.14117
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25=0.0042769
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25=0.00052637
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26=0.015878
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26=2.7094e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26=-3.8525e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26=-4782.4
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26=2.6665e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26=1.1346
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26=-0.0022969
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26=0.010965
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26=0.034452
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27=0.04327
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27=0.055573
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27=0.015383
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27=1.2388e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27=-1.4023e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27=-2900.8
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27=8.9139e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27=1.45
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27=-0.0047977
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28=6.9059e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28=1.5282
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28=-0.003291
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28=0.018194
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28=0.071288
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28=0.0074048
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28=-5.0866e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28=-1.027e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28=-0.00029663
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28=-3132.1
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29=6.6011e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29=2.3772
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29=-0.0019752
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29=0.076957
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29=0.11084
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29=-0.049364
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29=0.008623
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29=1.0863e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29=-4.4728e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29=-0.030186
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30=-0.019877
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30=6.7629e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30=3.0155
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30=-0.0011218
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30=0.098094
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30=0.0034884
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30=0.00077199
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30=1.0547e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30=-2.2772e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30=-0.00085806
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31=3.4884e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31=3.4223
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31=-0.002448
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31=0.021542
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31=0.12922
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31=0.0079843
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31=0.0029578
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31=1.463e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31=-5.4101e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31=0.0097768
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31=-0.0010532
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32=4.7775e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32=3.8903
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32=-0.0019471
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32=-0.21531
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32=0.16199
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32=0.0068898
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32=0.00046848
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32=1.0384e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32=-4.4536e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32=-0.0013947
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33=-4311.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33=2.4489e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33=1.3538
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33=-0.0030453
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33=-0.0073629
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33=0.036431
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33=0.019486
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33=2.8817e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33=-8.2061e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34=-2734.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34=1.4364e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34=1.6711
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34=-0.003633
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34=0.11006
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34=0.082979
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34=0.0080238
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34=3.887e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34=-1.0184e-18
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35=2.5095e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35=-0.0001809
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35=-0.032724
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35=6.1346e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35=1.2231e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35=9.0298e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35=1.7437
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35=0.00083875
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35=0.0066706
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35=0.060894
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35=0.0035595
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35=5.9894e-13
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36=4.7238e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36=8.7499e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36=2.3627e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36=1.0455e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36=4.5702e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36=4.444
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36=-5.5268e-5
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36=-0.64962
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36=0.14456
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36=-0.00025779
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37=-0.0013459
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37=-1.2717e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37=2.4827e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37=-0.044516
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37=6.7541e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37=6.4156e-8
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37=1.3311e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37=2.534
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37=0.0009913
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37=-0.22407
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37=0.073263
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38=-0.069099
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38=0.11229
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38=2.4551e-5
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38=3.9386e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38=2.2142e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38=0.0023234
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38=-0.040882
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38=6.659e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38=6.8754e-9
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38=8.2858e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38=3.7975
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38=0.00066016
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39=8.6355e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39=3.6502
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39=-0.00040288
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39=-0.16616
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39=0.14014
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39=0.0017461
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39=2.2233e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39=-6.3117e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39=0.0047338
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39=6.3852e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39=7.4391e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40=0.00075209
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40=3.6771e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40=0.44397
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40=-0.0042826
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40=0.13292
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40=0.031311
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40=-5.0918e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40=-1.8296e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40=-1.3739e-5
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40=-18056.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41=-0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41=0.022687
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41=7.191e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41=1.3473
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41=0.00015782
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41=0.093611
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41=0.013589
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41=-2.67e-13
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41=-8.3946e-20
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41=-0.00056891
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41=-11763.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42=-0.21909
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42=1.6489e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42=2.0237
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42=-0.0014079
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42=0.13849
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42=0.044229
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42=0.013318
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42=2.5227e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42=-1.1626e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42=-0.0036779
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42=-8835.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43=2.3794e-7
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43=2.867e-10
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43=5.9956e-10
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43=1.5498
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43=-0.0020643
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43=-0.033997
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43=0.095194
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43=0.0079272
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43=-2.503e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43=-8.6763e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43=0.00057915
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44=0.002216
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44=1.5134e-7
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44=3.504e-10
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44=8.9047e-10
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44=2.0398
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44=-0.0024078
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44=-0.1299
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44=0.10552
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44=0.0089111
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44=-2.2688e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44=-9.51e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45=0.0030097
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45=9.3768e-8
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45=3.0925e-10
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45=8.4822e-8
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45=3.5348
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45=-0.0012711
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45=-0.1231
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45=0.14185
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45=0.0053491
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45=-8.113e-14
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45=-3.3415e-19
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46=-1.3254e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46=-0.00191
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46=-10829.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46=4.3673e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46=0.36952
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46=-0.0034037
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46=0.065803
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46=0.083364
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46=0.023517
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46=-3.6609e-12
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47=-1.7538e-12
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47=-1.0172e-18
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47=-11219.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47=1.3897e-9
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47=1.8271
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47=-0.0030917
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47=0.053253
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47=0.10563
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47=0.011414
.param sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48=0.011228
.param sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48=-2.9549e-14
.param sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48=-1.2932e-19
.param sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48=-0.0010854
.param sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48=-8790.2
.param sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48=0.0
.param sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48=3.1236e-7
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48=1.3807
.param sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48=-0.00040428
.param sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48=0.036224
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48=0.066072
.include "sky130_fd_pr__pfet_g5v0d10v5.pm3.spice"