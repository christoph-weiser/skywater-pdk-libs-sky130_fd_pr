* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__nfet_05v0_nvt__toxe_mult=1.052
.param sky130_fd_pr__nfet_05v0_nvt__rshn_mult=1.0
.param sky130_fd_pr__nfet_05v0_nvt__overlap_mult=1.3700
.param sky130_fd_pr__nfet_05v0_nvt__ajunction_mult=1.3878e+0
.param sky130_fd_pr__nfet_05v0_nvt__pjunction_mult=1.2464e+0
.param sky130_fd_pr__nfet_05v0_nvt__lint_diff=-1.7325e-8
.param sky130_fd_pr__nfet_05v0_nvt__wint_diff=3.2175e-8
.param sky130_fd_pr__nfet_05v0_nvt__dlc_diff=-3.0000e-8
.param sky130_fd_pr__nfet_05v0_nvt__dwc_diff=3.2175e-8
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_0=-0.056577
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_0=0.08428
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_0=0.00016793
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_0=-0.005636
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_0=-1.9616e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_0=0.032906
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_0=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_0=0.0068039
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_0=-1.0516e-18
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_1=-1.0828e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_1=0.091002
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_1=0.042279
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_1=-0.0025266
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_1=-0.0056151
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_1=-2.4885e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_1=0.020743
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_1=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_1=0.004878
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_2=-1.0026e-18
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_2=-0.19806
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_2=0.0025007
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_2=-0.0058474
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_2=-1.9172e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_2=2871.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_2=0.040758
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_2=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_3=-1.2607e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_3=0.021014
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_3=-7.6708e-19
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_3=0.1208
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_3=0.00073216
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_3=-0.004008
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_3=-0.0057207
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_3=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_3=0.001698
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_4=-0.0061975
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_4=0.014978
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_4=-2.6745e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_4=0.033608
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_4=-1.0632e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_4=0.12546
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_4=0.1273
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_4=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_4=-0.001136
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_5=0.00076607
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_5=-0.0073364
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_5=0.012511
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_5=-1.8417e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_5=0.026896
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_5=-1.0258e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_5=0.12026
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_5=0.11694
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_5=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_6=0.062703
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_6=-0.0018694
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_6=-0.0057585
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_6=0.0066755
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_6=-1.5181e-11
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_6=0.013027
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_6=-8.6079e-19
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_6=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_6=0.15139
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_7=-0.062415
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_7=0.00069645
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_7=-0.0070762
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_7=0.020702
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_7=-2.2827e-11
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_7=3748.4
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_7=-1.0099e-18
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_7=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_8=0.010794
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_8=-2.5551e-8
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_8=0.0029018
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_8=-0.0068423
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_8=0.0021841
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_8=-6.2851e-12
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_8=3.5554e-10
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_8=-6.4524e-19
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_8=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_9=0.15402
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_9=0.004958
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_9=-0.0072966
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_9=0.035399
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_9=2.2764e-13
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_9=1592.8
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_9=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_9=-2.896e-19
.param sky130_fd_pr__nfet_05v0_nvt__vsat_diff_10=2509.5
.param sky130_fd_pr__nfet_05v0_nvt__vth0_diff_10=0.025399
.param sky130_fd_pr__nfet_05v0_nvt__b0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__keta_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__b1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__kt1_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pditsd_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__pclm_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__nfactor_diff_10=-0.019006
.param sky130_fd_pr__nfet_05v0_nvt__ags_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__u0_diff_10=-0.0078678
.param sky130_fd_pr__nfet_05v0_nvt__pdits_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__k2_diff_10=0.00080055
.param sky130_fd_pr__nfet_05v0_nvt__ua_diff_10=-1.5105e-11
.param sky130_fd_pr__nfet_05v0_nvt__eta0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__ub_diff_10=-7.9876e-19
.param sky130_fd_pr__nfet_05v0_nvt__tvoff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__voff_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__a0_diff_10=0.0
.param sky130_fd_pr__nfet_05v0_nvt__rdsw_diff_10=0.0
.include "sky130_fd_pr__nfet_05v0_nvt.pm3.spice"