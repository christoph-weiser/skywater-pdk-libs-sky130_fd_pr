* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.include "../../sonos_e/begin_of_life.pm3.spice"
.include "../../sonos_p/begin_of_life.pm3.spice"
.include "../../sonos_e/end_of_life/ff.spice"
.include "../../sonos_p/end_of_life/ff.spice"