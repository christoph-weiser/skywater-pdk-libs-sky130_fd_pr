* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__toxe_mult=1.06
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rbpb_mult=1.2
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__overlap_mult=1.0412
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__ajunction_mult=1.1726
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__pjunction_mult=1.2510
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__lint_diff=-1.7325e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__wint_diff=3.2175e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__rshg_diff=7.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dlc_diff=-1.7325e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_b__xgw_diff=6.4250e-8
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_0=0.061109
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_0=2277.3
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_0=0.0082757
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_0=-0.0032379
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vth0_diff_1=0.062761
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__vsat_diff_1=2408.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__k2_diff_1=0.01206
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__u0_diff_1=8.1975e-5
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_0=2239.7
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_0=0.051379
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_0=0.0080646
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_0=-0.0035332
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_1=-2.1067
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_1=0.055351
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_1=0.011508
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_1=-0.00040977
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vsat_diff_2=-617.15
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__vth0_diff_2=0.061066
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__k2_diff_2=0.0081582
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__u0_diff_2=-0.0027923
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_0=0.0074618
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_0=-0.0021786
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_0=0.061096
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_0=11951.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_1=0.0043804
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_1=-0.0025862
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_1=0.052501
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_1=-1288.1
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__k2_diff_2=0.0069032
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__pclm_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__u0_diff_2=-0.0090934
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vth0_diff_2=0.045939
.param sky130_fd_pr__rf_nfet_g5v0d10v5_bm10__vsat_diff_2=10578.0
.include "sky130_fd_pr__rf_nfet_g5v0d10v5_b.pm3.spice"