* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.param sky130_fd_pr__rf_nfet_01v8_b__toxe_mult=0.948
.param sky130_fd_pr__rf_nfet_01v8_b__rbpb_mult=0.8
.param sky130_fd_pr__rf_nfet_01v8_b__overlap_mult=0.94816
.param sky130_fd_pr__rf_nfet_01v8_b__ajunction_mult=0.7739
.param sky130_fd_pr__rf_nfet_01v8_b__pjunction_mult=0.79336
.param sky130_fd_pr__rf_nfet_01v8_b__lint_diff=1.7325e-8
.param sky130_fd_pr__rf_nfet_01v8_b__wint_diff=-3.2175e-8
.param sky130_fd_pr__rf_nfet_01v8_b__rshg_diff=-7.0
.param sky130_fd_pr__rf_nfet_01v8_b__dlc_diff=12.773e-9
.param sky130_fd_pr__rf_nfet_01v8_b__dwc_diff=0.0
.param sky130_fd_pr__rf_nfet_01v8_b__xgw_diff=-6.4250e-8
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_0=-0.075991
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_0=-22417.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_0=0.010085
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_0=0.00074749
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_1=-0.039487
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_1=-19233.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_1=0.020683
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_1=0.0011292
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_2=-0.043022
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_2=-16781.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_2=0.038033
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_2=0.0006468
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_3=-0.035105
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_3=-28463.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_3=0.010626
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_3=-0.0036794
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_4=-0.05182
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_4=-25171.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_4=0.030375
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_4=-0.0033229
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_5=-0.032322
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_5=-20257.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_5=0.042979
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_5=0.0011015
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_6=-0.0033456
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_6=-0.041439
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_6=-28660.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_6=0.0064952
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_7=0.02645
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_7=-0.0036669
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_7=-0.045761
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_7=-23039.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__k2_diff_8=0.04175
.param sky130_fd_pr__rf_nfet_01v8_bm02__u0_diff_8=-0.0010573
.param sky130_fd_pr__rf_nfet_01v8_bm02__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm02__vth0_diff_8=-0.032973
.param sky130_fd_pr__rf_nfet_01v8_bm02__vsat_diff_8=-16043.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_0=0.0091842
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_0=-0.00070926
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_0=-0.051501
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_0=-31984.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_0=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_1=0.028977
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_1=-0.0013648
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_1=-0.058125
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_1=-23564.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_1=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_2=0.042169
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_2=-0.00035031
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_2=-0.046633
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_2=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_2=-19030.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_3=-30928.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_3=0.013856
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_3=-0.0048131
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_3=-0.046817
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_3=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_4=-24921.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_4=0.034977
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_4=-0.0071423
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_4=-0.061148
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_4=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_5=-8528.2
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_5=0.045401
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_5=-0.0043436
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_5=-0.04118
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_5=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_6=-29958.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_6=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_6=0.009601
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_6=-0.0033405
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_6=-0.04502
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_7=-0.0060347
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_7=-26996.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_7=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_7=0.031931
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_7=-0.060436
.param sky130_fd_pr__rf_nfet_01v8_bm04__vth0_diff_8=-0.0389
.param sky130_fd_pr__rf_nfet_01v8_bm04__u0_diff_8=-0.0030982
.param sky130_fd_pr__rf_nfet_01v8_bm04__b1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__voff_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__kt1_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ub_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__nfactor_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__vsat_diff_8=-11896.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ags_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__a0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__b0_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__ua_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__rdsw_diff_8=0.0
.param sky130_fd_pr__rf_nfet_01v8_bm04__k2_diff_8=0.044114
.include "sky130_fd_pr__rf_nfet_01v8_b.pm3.spice"